@00000000
18000000
A8200001
C0000811
C1400000
18800000
A8840120
44002000
15000000
04000254
15000000
04000002
15000000
15000000
00000002
15000000
9C200001
9C410002
9C620004
9C830008
9CA40010
9CC50020
9CE60040
9D070080
9D280100
9D490200
9D6A0400
9D8B0800
9DAC1000
9DCD2000
9DEE4000
9E0F8000
E3E00802
E3DF1002
E3BE1802
E39D2002
E37C2802
E35B3002
E33A3802
E3194002
E2F84802
E2D75002
E2B65802
E2956002
E2746802
E2537002
E2327802
E2118002
1BE00000
ABFF0040
C0408234
D41F8000
18601234
A8635678
D41F1804
8C9F0004
E1082000
D81F200B
8C9F0005
E1082000
D81F200A
8C9F0006
E1082000
D81F2009
8C9F0007
E1082000
D81F2008
909F0008
E1082000
D81F2007
909F0009
E1082000
D81F2006
909F000A
E1082000
D81F2005
909F000B
E1082000
D81F2004
949F0004
E1082000
DC1F200A
949F0006
E1082000
DC1F2008
989F0008
E1082000
DC1F2006
989F000A
E1082000
DC1F2004
849F0004
E1082000
C0404234
853F0000
E1094000
D41F4000
9C600001
9C800002
9CA0FFFF
9CC0FFFF
9D000000
E0E51802
E1032802
E1083800
E1232000
E0E93B06
E1083800
C0404234
853F0000
E1094000
D41F4000
9C600001
9C800002
9CA0FFFF
9CC0FFFF
9D000000
A5080001
E1081803
AD05A5A5
E1082805
A9080002
E1082004
C0404234
853F0000
E1094000
D41F4000
9C600001
9C800002
9CA0FFFF
9CC0FFFF
9D000000
B9050006
E1082008
B9080046
E1082048
B9080082
E1082088
C0404234
853F0000
E1094000
D41F4000
9C600001
9C80FFFE
9D000000
E4031800
B4A00011
A4850200
E1082000
E4032000
B4A00011
A4850200
E1082000
BC030001
B4A00011
A4850200
E1082000
BC03FFFE
B4A00011
A4850200
E1082000
E4231800
B4A00011
A4850200
E1082000
E4232000
B4A00011
A4850200
E1082000
BC230001
B4A00011
A4850200
E1082000
BC23FFFE
B4A00011
A4850200
E1082000
E4431800
B4A00011
A4850200
E1082000
E4432000
B4A00011
A4850200
E1082000
BC430001
B4A00011
A4850200
E1082000
BC43FFFE
B4A00011
A4850200
E1082000
E4631800
B4A00011
A4850200
E1082000
E4632000
B4A00011
A4850200
E1082000
BC630001
B4A00011
A4850200
E1082000
BC63FFFE
B4A00011
A4850200
E1082000
E4831800
B4A00011
A4850200
E1082000
E4832000
B4A00011
A4850200
E1082000
BC830001
B4A00011
A4850200
E1082000
BC83FFFE
B4A00011
A4850200
E1082000
E4A31800
B4A00011
A4850200
E1082000
E4A32000
B4A00011
A4850200
E1082000
BCA30001
B4A00011
A4850200
E1082000
BCA3FFFE
B4A00011
A4850200
E1082000
E5431800
B4A00011
A4850200
E1082000
E5432000
B4A00011
A4850200
E1082000
BD430001
B4A00011
A4850200
E1082000
BD43FFFE
B4A00011
A4850200
E1082000
E5631800
B4A00011
A4850200
E1082000
E5632000
B4A00011
A4850200
E1082000
BD630001
B4A00011
A4850200
E1082000
BD63FFFE
B4A00011
A4850200
E1082000
E5831800
B4A00011
A4850200
E1082000
E5832000
B4A00011
A4850200
E1082000
BD830001
B4A00011
A4850200
E1082000
BD83FFFE
B4A00011
A4850200
E1082000
E5A31800
B4A00011
A4850200
E1082000
E5A32000
B4A00011
A4850200
E1082000
BDA30001
B4A00011
A4850200
E1082000
BDA3FFFE
B4A00011
A4850200
E1082000
C0404234
853F0000
E1094000
D41F4000
9DC00004
9DE00014
9EA00040
9E000010
9E200007
9E400008
9E600009
9E80FFFF
D40E0000
D40E0004
D40E0008
D40E000C
D40E0010
D40E0014
D40E0018
D40E001C
D40E0020
D40E0024
D40E0028
D40E002C
9DC00004
9E000010
E2317000
E2319800
E231A005
9E10FFFC
9DCE0004
BC100000
10000004
E2319000
03FFFFF8
9E730001
9DC00004
9E000010
E2317000
E2319800
E231A005
9E10FFFC
9DCE0004
E46E7800
10000004
E2319000
03FFFFF8
9E710001
9DC00004
9E000010
E2317000
E2319800
E231A005
9E10FFFC
9DCE0004
BC100000
10000004
E2317000
03FFFFF8
B2730002
9DC00004
9E000010
E2317000
E2319800
E231A005
9E10FFFC
9DCE0004
E46E7800
10000004
E2317000
03FFFFF8
B2710001
9DC00004
9E000010
E2317000
E2319800
E231A005
9E10FFFC
9DCE0004
BC100000
10000004
E2319306
03FFFFF8
9E730001
9DC00004
9E000010
E2317000
E2319800
E231A005
9E10FFFC
9DCE0004
E46E7800
10000004
E2319306
03FFFFF8
9E710001
9DC00004
9E000010
E2317000
E2319800
E231A005
9E10FFFC
9DCE0004
BC100000
10000004
E2317306
03FFFFF8
B2730002
9DC00004
9E000010
E2317000
E2319800
E231A005
9E10FFFC
9DCE0004
E46E7800
10000004
E2317306
03FFFFF8
B2710001
9DC00004
9E000010
E2317000
E2319800
E231A005
9E10FFFC
B1CE0002
BC100000
10000004
E2319000
03FFFFF8
9E730001
9DC00004
9E000010
E2317000
E2319800
E231A005
9E10FFFC
B1CE0002
E46EA800
10000004
E2319000
03FFFFF8
9E710001
9DC00004
9E000010
E2317000
E2319800
E231A005
9E10FFFC
B1CE0002
BC100000
10000004
E2317000
03FFFFF8
B2730002
9DC00004
9E000010
E2317000
E2319800
E231A005
9E10FFFC
B1CE0002
E46EA800
10000004
E2317000
03FFFFF8
B2710001
9DC00004
9E000010
E2317000
E2319800
E231A005
9E10FFFC
B1CE0002
BC100000
10000004
E2319306
03FFFFF8
9E730001
9DC00004
9E000010
E2317000
E2319800
E231A005
9E10FFFC
B1CE0002
E46EA800
10000004
E2319306
03FFFFF8
9E710001
9DC00004
9E000010
E2317000
E2319800
E231A005
9E10FFFC
B1CE0002
BC100000
10000004
E2317306
03FFFFF8
B2730002
9DC00004
9E000010
E2317000
E2319800
E231A005
9E10FFFC
B1CE0002
E46EA800
10000004
E2317306
03FFFFF8
B2710001
9DC00004
9E000010
E2317000
E231A005
9E10FFFC
9DCE0004
E46E7800
0FFFFFFB
D4108800
9DC00004
9E000010
E231B000
E2317000
E231A005
9E10FFFC
9DCE0004
E46E7800
0FFFFFFA
86D00000
E231B000
E231A005
04000006
B2310002
E2319000
E231A005
00000006
E2528802
9E310001
E231A005
44004800
9E520008
E2319306
1A40B093
AA52A787
E2319002
15000000
15000000
E1008800
00000005
9D080001
E1404804
48005000
9D080001
07FFFFFD
9D080001
BC000000
10000002
9D080001
BC000001
10000003
9D080001
9D080001
BC000000
0C000003
9D080001
9D080001
BC000001
0C000003
9D080001
9D080001
18600000
A8630A30
C0001820
B4A00011
C0002840
24000000
9D080001
9D080001
C0404234
853F0000
E1094000
D41F4000
853F0000
1860CC69
A863E5FB
E0681800
18805EAD
A884DEA0
E0632002
15000002
A8600000
15000001
15000000
15000000
B4600001
A4830004
E4040000
10000021
15000000
B4C00011
9CA0FFFF
ACA50010
E0A62803
C0002811
B4600006
A4830080
B8A40047
A8C00010
E1C62808
A4830078
B8A40043
A8C00001
E0E62808
9CC00000
E0AE2808
C0803002
E4262800
13FFFFFE
E0C67000
B4C00011
A8C60010
C0003011
15000000
15000000
15000000
15000000
15000000
15000000
15000000
15000000
B4600001
A4830002
E4040000
10000019
15000000
B4C00011
9CA0FFFF
ACA50008
E0A62803
C0002811
B4600005
A4830080
B8A40047
A8C00010
E1C62808
A4830078
B8A40043
A8C00001
E0E62808
9CC00000
E0AE2808
C0603003
E4262800
13FFFFFE
E0C67000
B4C00011
A8C60008
C0003011
44004800
15000000
	 
