@00000000
18000000
18A0FFFF
A8A5FFFF
E0C50004
18809100
A8842000
D4042804
D4043000
E0C62805
18E00010
9CE7FFFF
E4070000
0FFFFFFE
15000000
03FFFFF9
15000000
	 
