@00000000
18000000
04000018
15000000
04000040
15000000
0400005B
15000000
15000002
15000001
E1630000
15000000
04000040
15000000
B8E30008
04000052
15000000
E0E71800
E0670004
15000000
15000001
15000000
A860DEAD
15000002
15000001
15000000
18809000
A8840000
9CA00080
D8042803
9CA00024
D8042800
9CA00000
D8042801
9CA00003
D8042803
9CA000C3
D8042802
9CA00000
D8042801
44004800
15000000
19009000
A9080000
8C680005
A4630001
BC030000
13FFFFFD
15000000
8C680000
44004800
15000000
04000018
B8830010
04000016
B8A30018
E0C42804
44004800
15000000
E0863800
18A00000
0400000F
E1442800
9CA50001
D80A1800
E4055000
0FFFFFFB
15000000
E1890004
07FFFFE5
15000000
BC03003A
0FFFFFFD
15000000
44006000
15000000
E1890004
07FFFFDD
15000000
BCA30030
13FFFFC6
15000000
BC830039
0C000005
15000000
9C63FFD0
44006000
15000000
BCA30041
13FFFFBD
15000000
BCA30046
0FFFFFBA
15000000
9C63FFC9
44006000
15000000
E1A90004
07FFFFEA
15000000
B9C30004
07FFFFE7
15000000
E06E1804
44006800
15000000
	 
