@00000000
18000000
18400000
18A00000
18C00000
A8C60100
18E00000
18400102
A8420304
D4071000
84270000
18401819
A8421A1B
D4071004
84270004
18402829
A8422A2B
D4071008
84270008
18403839
A8423A3B
D407100C
8427000C
18404849
A8424A4B
D4071010
84270010
18405859
A8425A5B
D4071014
84270014
18406869
A8426A6B
D4071018
84270018
18407879
A8427A7B
D407101C
8427001C
18408889
A8428A8B
D4071020
84270020
18409899
A8429A9B
D4071024
84270024
1840A8A9
A842AAAB
D4071028
84270028
1840B8B9
A842BABB
D407102C
8427002C
18E00100
18401112
A8421314
D4071000
84270000
18E00200
18402122
A8422324
D4071000
84270000
18E00300
18403132
A8423334
D4071000
84270000
18E00400
18404142
A8424344
D4071000
84270000
18E00500
18405152
A8425354
D4071000
84270000
18E00600
18406162
A8426364
D4071000
84270000
18E00700
18407172
A8427374
D4071000
84270000
18E09600
A8E70000
18400000
A842FFFF
D4071008
18400000
18809100
A8840000
D4040004
84A40000
A4A52000
BC050000
13FFFFFD
15000000
44003000
15000000
	 
