@00000000
18000000
18200000
18400000
18600000
18800000
18A00000
18C00000
18E00000
19000000
19200000
19400000
19600000
19800000
19A00000
19C00000
19E00000
1A000000
1A200000
1A400000
1A600000
1A800000
1AA00000
1AC00000
1AE00000
1B000000
1B200000
1B400000
1B600000
1B800000
1BA00000
1BC00000
1BE00000
A8200001
C0000811
C1400000
18800000
A8842030
44002000
15000000
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
000017BF
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
0000177F
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
0000173F
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
000016FF
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
000016BF
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
0000167F
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
0000163F
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
000015FF
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
000015BF
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
0000157F
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
0000153F
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
000014FF
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
000014BF
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
0000147F
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
0000143F
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
000013FF
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
000013BF
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
0000137F
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
0000133F
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
000012FF
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
000012BF
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
0000127F
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
0000123F
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
000011FF
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
000011BF
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
0000117F
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
0000113F
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
000010FF
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
000010BF
B4800020
D4000804
18200000
A8219C0C
84210000
E4010000
0C000006
15000000
18200000
A8219C10
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600000
A8639C0C
84830000
9C840001
D4032000
B4600010
0000107F
B4800020
15000000
15000000
9C21FFFC
D4014800
040000BC
15000000
04001351
15000000
85210000
44004800
9C210004
44004800
15000000
04000FE3
15000000
040012E4
15000000
18600000
A8639A8C
18800000
A8849C98
D4030000
E4832000
13FFFFFE
9C630004
18200000
A8216BA4
84210000
18400000
A8426BA8
84420000
E0211000
18600000
A8639C10
D4030800
18600000
A8638E1C
84630000
E0811802
18A00000
A8A59C18
D4052000
E0202004
E0410804
18600000
A8639C14
D4030800
18600000
A8638E18
84630000
E0811802
18A00000
A8A59C1C
D4052000
0400118A
15000000
0400111D
15000000
07FFFFC8
15000000
18600000
040000BB
A8636DC8
18800000
A8846BB0
84840000
E4240000
0C000004
E0600004
04000F3E
15000000
040012AE
15000000
E0600004
E0800004
0400009C
E0A00004
040000B7
9C6B0000
15000000
D7E117F8
18600000
18400000
A8639A8F
A8429A8C
D7E14FFC
E0631002
D7E10FF4
BCA30006
10000009
9C21FFF4
18800000
A8840000
BC040000
10000004
15000000
48002000
A8620000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E117F8
18600000
18400000
A8639A8C
A8429A8C
D7E14FFC
E0631002
D7E10FF4
B8630082
B883005F
E0841800
B8840081
BC040000
10000009
9C21FFF4
18A00000
A8A50000
BC050000
10000004
15000000
48002800
A8620000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E197F8
1A400000
D7E117F0
AA529A8C
D7E14FFC
8C520000
D7E10FEC
D7E177F4
BC220000
10000026
9C21FFEC
19C00000
18800000
A9CE8E10
A8848E0C
18400000
E1CE2002
A8429A90
B9CE0082
84620000
9DCEFFFF
E4837000
0C00000E
9C630001
18A00000
B8830002
A8A58E0C
D4021800
E0642800
84630000
48001800
15000000
84620000
E4837000
13FFFFF6
9C630001
07FFFFAA
18400000
A8420000
BC220000
0C000006
9C400001
18600000
07FFF753
A8638E00
9C400001
D8121000
9C210014
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
D7E14FFC
D7E10FF8
9C21FFF8
9C210008
8521FFFC
44004800
8421FFF8
18600000
D7E14FFC
A8630000
D7E10FF8
BC030000
10000007
9C21FFF8
18600000
18800000
A8638E00
07FFF737
A8849A94
18600000
A8638E14
84830000
BC040000
0C000008
18800000
07FFFF96
15000000
9C210008
8521FFFC
44004800
8421FFF8
A8840000
BC040000
13FFFFF8
15000000
48002000
15000000
03FFFFF4
15000000
D7E14FFC
D7E10FF8
9C21FFF8
9C210008
8521FFFC
44004800
8421FFF8
D7E117F8
9C410000
D7E14FFC
9C21FFF0
D7E21FF4
D7E227F0
18600000
A8636DE4
0400005D
15000000
9C600000
A9630000
A8220000
8441FFF8
8521FFFC
44004800
15000000
A8830000
9C600000
D7E14FFC
D7E10FF8
A8A30000
9C21FFF8
0400009E
A8C30000
9C210008
8521FFFC
44004800
8421FFF8
D7E117F8
D7E14FFC
D7E10FF4
9C800000
9C21FFF4
040000E3
A8430000
18600000
A8636DF4
84630000
8483003C
BC040000
10000004
15000000
48002000
15000000
04000DE1
A8620000
D7E117F4
D7E177F8
A8440000
A9C30000
D7E14FFC
A8640000
D7E10FF0
0400003D
9C21FFD4
D401100C
18400000
9C8B0001
A8426DFA
846E0038
D4011014
9C400001
D4015810
D4011018
9C41000C
D4012008
D4011000
9C400002
BC230000
D4011004
0C00001A
844E0008
9862000C
A4832000
BC240000
10000007
9CA0DFFF
84820064
A8632000
E0842803
DC02180C
D4022064
A86E0000
A8820000
0400025F
A8A10000
BC2B0000
10000003
9D60FFFF
9D60000A
9C21002C
8521FFFC
8421FFF0
8441FFF4
44004800
85C1FFF8
0400021B
A86E0000
03FFFFE7
9862000C
D7E14FFC
D7E117F8
D7E10FF4
9C21FFF4
04000427
A8430000
A8820000
07FFFFC3
A86B0000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
A4830003
D7E10FF8
D7E117FC
BC040000
1000003A
9C21FFF8
90A30000
BC050000
10000038
A8830000
00000007
9C840001
90A40000
BC250000
0C00002C
E1641802
9C840001
A4A40003
BC250000
13FFFFF9
15000000
1840FEFE
84A40000
A842FEFF
E0C51000
ACA5FFFF
18408080
E0A62803
A8428080
E0A51003
BC250000
10000010
15000000
9C840004
1840FEFE
84A40000
A842FEFF
E0C51000
ACA5FFFF
18408080
E0A62803
A8428080
E0A51003
BC050000
13FFFFF6
9C840004
9C84FFFC
90A40000
BC050000
10000009
E1641802
9C840001
90A40000
BC250000
13FFFFFE
9C840001
9C84FFFF
E1641802
9C210008
8421FFF8
44004800
8441FFFC
03FFFFD7
A8830000
03FFFFFA
A9650000
D7E117E8
18400000
D7E177EC
A8426DF4
D7E197F0
85C20000
D7E1A7F4
850E0148
D7E1B7F8
D7E14FFC
D7E10FE4
BC280000
9C21FFE4
AAC30000
A8440000
AA850000
0C00003B
AA460000
84E80004
BD47001F
10000014
18600000
BC360000
10000025
9CA70001
9CE70002
D4082804
B8E70002
9D600000
E0E83800
D4071000
9C21001C
8521FFFC
8421FFE4
8441FFE8
85C1FFEC
8641FFF0
8681FFF4
44004800
86C1FFF8
A8630000
BC230000
0FFFFFF5
9D60FFFF
07FFF639
9C600190
BC0B0000
1000001F
A90B0000
846E0148
9C800000
D40B1800
D40B2004
D40E5948
D40B2188
D40B218C
BC360000
9CA00001
0FFFFFDF
A8E40000
B9670002
9C800001
BC360002
E0685800
E0843808
D403A088
84C80188
E0C62004
D4083188
13FFFFD4
D4039108
8468018C
E0832004
03FFFFD0
D408218C
9D0E014C
03FFFFC6
D40E4148
03FFFFD1
9D60FFFF
D7E117D8
18400000
D7E1F7F8
A8426DF4
D7E197E0
87C20000
D7E1D7F0
D7E1E7F4
D7E14FFC
D7E10FD4
D7E177DC
D7E1A7E4
D7E1B7E8
D7E1C7EC
9C5E0148
9C21FFD0
1B800000
AB430000
AA440000
D4011000
AB9C0000
869E0148
BC340000
0C000043
86C10000
84540004
9DC2FFFF
BD6E0000
0C00002F
BC1C0000
9C420001
B8420002
0000000A
E0541000
84620100
E4039000
10000009
15000000
9DCEFFFF
BC2EFFFF
0C000022
9C42FFFC
BC120000
0FFFFFF7
15000000
84740004
9C63FFFF
E4237000
0C000041
84A20000
9C600000
D4021800
BC050000
13FFFFF1
9C600001
E0837008
84740188
E0641803
BC030000
0C00002C
87140004
48002800
15000000
84740004
E423C000
13FFFFD4
15000000
84760000
E423A000
13FFFFD0
9DCEFFFF
BC2EFFFF
13FFFFE2
9C42FFFC
BC1C0000
1000000F
15000000
84540004
BC220000
10000028
84540000
BC020000
10000025
A8740000
07FFF5C1
D4161000
86960000
BC340000
13FFFFC1
15000000
9C210030
8521FFFC
8421FFD4
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
8474018C
E0641803
BC230000
10000009
15000000
A87A0000
48002800
84820080
03FFFFD1
84740004
03FFFFC3
D4147004
48002800
84620080
03FFFFCB
84740004
AAD40000
03FFFFDF
AA820000
D7E10FFC
9C21FFFC
9D600000
9C210004
44004800
8421FFFC
D7E10FFC
9C21FFFC
9D600000
9C210004
44004800
8421FFFC
18800000
D7E14FFC
D7E10FF8
A8844F34
040002CC
9C21FFF8
9C210008
8521FFFC
44004800
8421FFF8
18800000
D7E1A7E4
A88429C4
AA830000
D7E14FFC
D7E117D8
D7E177DC
D7E197E0
D7E1B7E8
D7E1C7EC
D7E1D7F0
D7E1E7F4
D7E1F7F8
D7E10FD4
9C400000
D414203C
9C6302EC
9C800003
85D40004
9CC00004
D41412E0
D41422E4
D4141AE8
9C21FFD4
9C6E005C
A8820000
D40E1000
D40E1004
D40E1008
DC0E300C
D40E1064
DC0E100E
D40E1010
D40E1014
D40E1018
9CA00008
1B800000
1B400000
1B000000
0400064D
1AC00000
AB9C4BE0
AB5A4C60
AB184CF0
AAD64D58
86540008
9FC00001
9CC00009
D40EE020
D40ED024
D40EC028
D40EB02C
D40E701C
9C72005C
A8820000
D4121000
D4121004
D4121008
DC12300C
D4121064
DC12F00E
D4121010
D4121014
D4121018
04000634
9CA00008
9C600012
85D4000C
9CC00002
D412E020
D412D024
D412C028
D412B02C
D412901C
D40E1000
D40E1004
D40E1008
DC0E180C
D40E1064
D40E1010
D40E1014
D40E1018
DC0E300E
9C6E005C
A8820000
0400061F
9CA00008
D40EE020
D40ED024
D40EC028
D40EB02C
D40E701C
D414F038
9C21002C
8521FFFC
8421FFD4
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
D7E117F0
D7E177F4
9C44FFFF
9DC00068
D7E197F8
E1C27306
D7E14FFC
D7E10FEC
AA440000
9C21FFEC
04000289
9C8E0074
BC0B0000
10000009
A84B0000
9C6B000C
9C800000
D40B9004
D40B2000
D40B1808
040005F6
9CAE0068
9C210014
A9620000
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
D7E117F0
18400000
D7E177F4
A8426DF4
D7E197F8
85C20000
D7E14FFC
844E0038
D7E10FEC
BC220000
9C21FFEC
10000004
AA430000
07FFFF6B
A86E0000
9DCE02E0
84AE0004
9CA5FFFF
BD850000
10000011
844E0008
9862000C
BC030000
10000013
9C820074
00000007
9CA5FFFF
98C4FF98
BC060000
1000000E
9C60FFFF
9CA5FFFF
9C44FFF4
BC25FFFF
13FFFFF9
9C840068
844E0000
BC220000
0C000021
15000000
03FFFFE8
A9C20000
9C60FFFF
9C800000
DC02180E
9C600001
9CA00008
DC02180C
9C600000
D4021864
D4021800
D4021808
D4021804
D4021810
D4021814
D4021818
040005B4
9C62005C
9C600000
A9620000
D4021830
D4021834
D4021844
D4021848
9C210014
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
A8720000
07FFFF9A
9C800004
BC0B0000
10000004
D40E5800
03FFFFC3
A9CB0000
9C40000C
03FFFFF0
D4121000
18600000
18800000
A8636DF4
D7E14FFC
D7E10FF8
A8844F34
9C21FFF8
040001E5
84630000
9C210008
8521FFFC
44004800
8421FFF8
84830038
D7E14FFC
D7E10FF8
BC240000
10000004
9C21FFF8
07FFFF13
15000000
9C210008
8521FFFC
44004800
8421FFF8
D7E10FFC
9C21FFFC
9C210004
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C210004
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C210004
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C210004
44004800
8421FFFC
D7E14FFC
D7E10FF8
040001F2
9C21FFF8
18800000
A86B0000
04000183
A8842994
9C210008
8521FFFC
44004800
8421FFF8
D7E14FFC
D7E10FF8
040001E6
9C21FFF8
18800000
A86B0000
04000177
A88429AC
9C210008
8521FFFC
44004800
8421FFF8
84C50008
D7E14FFC
D7E10FD4
D7E117D8
D7E177DC
D7E197E0
D7E1A7E4
D7E1B7E8
D7E1C7EC
D7E1D7F0
D7E1E7F4
D7E1F7F8
BC260000
0C00002C
9C21FFCC
94C4000C
ABC30000
A4660008
A8440000
BC030000
10000033
AA850000
84640010
BC230000
0C00002F
A6460002
A652FFFF
BC120000
10000037
85D40000
9EC00000
1B007FFF
AA560000
AB18FC00
BC120000
A8B60000
A87E0000
10000074
A8D20000
18807FFF
A884FC00
E4B22000
10000003
8482001C
A8D80000
85620024
48005800
15000000
BDAB0000
1000007F
E2D65800
84740008
E2525802
E1635802
BC2B0000
13FFFFEB
D4145808
9D600000
9C210034
8521FFFC
8421FFD4
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
A87E0000
0400077D
A8820000
BC2B0000
10000120
15000000
94C2000C
A6460002
A652FFFF
BC120000
0FFFFFCD
85D40000
A6C60001
BC160000
10000060
AB920000
D4019000
AAD20000
BC160000
1000003A
9C600000
84810000
BC240000
0C0000B7
A87C0000
E4B2B000
10000003
AB120000
AB160000
84C20014
84620008
AB580000
E0661800
D4011804
84620000
84810004
E5582000
10000003
9C800001
9C800000
A48400FF
BC040000
1000000B
E5983000
84A20010
E4432800
10000003
9C800001
9C800000
A48400FF
BC040000
0C0000D0
E5983000
10000082
A89C0000
85620024
A87E0000
8482001C
48005800
A8BC0000
BD4B0000
0C00002C
AB4B0000
E252D002
BC320000
0C000082
A87E0000
84740008
E39CD000
E063D002
E2D6D002
BC230000
0FFFFFAA
D4141808
BC160000
0FFFFFCA
9C600000
878E0000
86CE0004
D4011800
03FFFFC2
9DCE0008
86CE0000
864E0004
03FFFF87
9DCE0008
18607FFF
A863FFFF
E4B21800
10000005
A8720000
18800000
A8846DFC
84640000
04000EFE
A8980000
E0D85B06
A87E0000
85620024
8482001C
48005800
A8B60000
BD4B0000
10000021
15000000
9862000C
A8630040
9D60FFFF
03FFFF87
DC02180C
AA560000
BC120000
10000022
15000000
A4660200
BC030000
10000022
87820008
E492E000
10000053
AB1C0000
A4660480
BC230000
1000005D
15000000
84620000
A8960000
04000426
A8B80000
84620008
84820000
E383E002
E304C000
D402E008
D402C000
A9720000
84740008
E2D65800
E0635802
E2525802
BC030000
13FFFF65
D4141808
BC120000
0FFFFFE2
94C2000C
86CE0000
864E0004
03FFFFDB
9DCE0008
84620000
84820010
E4432000
10000006
E4B2E000
87020014
E472C000
13FFFFB9
E4B2E000
10000003
AB120000
AB1C0000
A8960000
04000402
A8B80000
84620008
84820000
E063C002
E084C000
D4021808
BC030000
10000004
D4022000
03FFFFDB
A9780000
A87E0000
04000869
A8820000
BC2B0000
13FFFFB6
15000000
03FFFFD3
A9780000
A8B80000
040003ED
E252D002
84620008
84820000
E063C002
E304C000
D4021808
BC320000
13FFFF83
D402C000
A87E0000
04000856
A8820000
BC0B0000
0FFFFFA3
15000000
03FFFF7B
D4019000
AB920000
84620000
03FFFFB2
AB120000
9C80000A
0400032A
A8B60000
BC0B0000
1000004E
9D6B0001
9C600001
E24BE002
03FFFF43
D4011800
84620014
84820010
E3031800
87420000
E0781800
E35A2002
BB03005F
9CFA0001
E0781800
E0E79000
BB030081
E4783800
10000004
A8B80000
AB070000
A8A70000
A4C60400
BC060000
10000028
A87E0000
040000AB
A8850000
BC2B0000
0C000037
AB8B0000
A86B0000
84820010
0400035B
A8BA0000
9462000C
9C80FB7F
E0632003
A8630080
DC02180C
E07CD000
E358D002
D402E010
D402C014
D4021800
AB920000
D402D008
03FFFF7D
AB120000
A89C0000
040003A1
84A10004
84A20000
84810004
A87E0000
E0A52000
A8820000
0400080E
D4022800
BC0B0000
0FFFFF5B
87410004
03FFFF30
E252D002
04000497
15000000
BC2B0000
13FFFFE5
AB8B0000
A87E0000
0400088E
84820010
9862000C
9C80FF7F
E0632003
9C80000C
03FFFF4C
D41E2000
9C800001
9E560001
03FFFEF7
D4012000
03FFFECF
9D60FFFF
9C80000C
9862000C
03FFFF42
D41E2000
D7E1B7F4
9EC302E0
D7E14FFC
D7E10FE0
D7E117E4
D7E177E8
D7E197EC
D7E1A7F0
D7E1C7F8
BC160000
1000002A
9C21FFE0
AB040000
9E800000
85D60004
9DCEFFFF
BD8E0000
10000014
86560008
9C52000C
9E52000E
94A20000
BCA50001
9DCEFFFF
10000009
9C62FFF4
98920000
BC04FFFF
10000006
BC2EFFFF
4800C000
15000000
E2945804
BC2EFFFF
9C420068
13FFFFF2
9E520068
86D60000
BC360000
13FFFFE7
15000000
9C210020
A9740000
8521FFFC
8421FFE0
8441FFE4
85C1FFE8
8641FFEC
8681FFF0
86C1FFF4
44004800
8701FFF8
03FFFFF5
AA960000
D7E1B7F4
9EC302E0
D7E14FFC
D7E10FE0
D7E117E4
D7E177E8
D7E197EC
D7E1A7F0
D7E1C7F8
BC160000
10000029
9C21FFE0
AB040000
AA830000
9E400000
85D60004
9DCEFFFF
BD8E0000
10000012
84560008
9C42000C
94A20000
BCA50001
9DCEFFFF
10000009
9C82FFF4
98A20002
BC05FFFF
10000005
A8740000
4800C000
15000000
E2525804
BC2EFFFF
13FFFFF3
9C420068
86D60000
BC360000
13FFFFE9
15000000
9C210020
A9720000
8521FFFC
8421FFE0
8441FFE4
85C1FFE8
8641FFEC
8681FFF0
86C1FFF4
44004800
8701FFF8
03FFFFF5
AA560000
00000C3C
15000000
D7E177DC
9DC4000B
D7E197E0
D7E14FFC
D7E10FD4
D7E117D8
D7E1A7E4
D7E1B7E8
D7E1C7EC
D7E1D7F0
D7E1E7F4
D7E1F7F8
BCAE0016
9C21FFD0
10000035
AA430000
9C40FFF8
E1CE1003
B86E005F
BC230000
10000036
E4447000
10000003
9C400001
A8430000
A44200FF
BC020000
0C000030
9C40000C
040003B4
A8720000
BC4E01F7
1000002E
18800000
A8849254
E06E2000
8443000C
E4221800
0C00015F
B8AE0043
84820004
9CA0FFFC
8462000C
E0842803
84C20008
E0822000
D406180C
84A40004
D4033008
A8A50001
A8720000
040003C8
D4042804
9D620008
9C210030
8521FFFC
8421FFD4
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
BC440010
10000007
9C40000C
0400038B
9DC00010
03FFFFDA
18800000
9C40000C
9D600000
03FFFFEA
D4121000
B8AE0049
BC050000
1000008A
BC450004
100000BD
BC450014
B8AE0046
9CC50038
E0A63000
18E00000
B8A50002
A8E79254
E0A53800
8445000C
E4051000
10000019
9D60FFFC
84620004
E0635803
E0837002
BD44000F
1000007A
BD640000
0C00000D
15000000
00000079
E0621800
9C80FFFC
84620004
E0632003
E0837002
BDA4000F
0C00006F
BD840000
0C00006F
15000000
8442000C
E4251000
13FFFFF5
15000000
9CA60001
1A800000
AA949254
84540010
9D140008
E4224000
0C000107
9CC0FFFC
84620004
E0633003
E0837002
BDA4000F
0C0000F2
BD840000
D4144014
0C000066
D4144010
BC4301FF
10000090
B8830049
B8630043
9CE00001
84940004
E0C31800
B8630082
B8C60002
E0671808
18E00000
A8E79254
E0632004
E0C63800
D4141804
84E60008
D402300C
D4023808
D4061008
D407100C
B8450082
9CC00001
E0C61008
E4461800
10000054
E0433003
BC220000
1000000F
E1652800
9C40FFFC
E0C63000
E0A51003
E0433003
BC220000
10000007
9CA50004
E0C63000
E0433003
BC020000
13FFFFFD
9CA50004
E1652800
18600000
B96B0002
A8639254
A9A50000
E16B1800
9D8B000C
9CECFFF4
844C0000
E4023800
10000019
9C80FFFC
84620004
E0632003
E0837002
BD44000F
100000CC
BD640000
0C00000D
E0821800
000000D2
84C2000C
9C80FFFC
84620004
E0632003
E0837002
BDA4000F
0C0000C1
BD840000
0C0000C7
15000000
8442000C
E4223800
13FFFFF5
15000000
9DAD0001
A44D0003
BC220000
13FFFFE1
9D8C0008
000000D5
A4650003
9CA0007E
03FFFF7C
9CC0003F
03FFFF99
9CC6FFFF
E0621800
84A2000C
84830004
84C20008
A8840001
D406280C
D4053008
D4032004
04000314
A8720000
03FFFF4D
9D620008
E0821800
A8720000
84A40004
A8A50001
0400030C
D4042804
03FFFF45
9D620008
84540008
9CA0FFFC
87020004
E3182803
E0787002
BDA3000F
10000003
9C800001
9C800000
A48400FF
BC240000
1000003A
E4987000
0C0000A2
9CA00001
A4A500FF
BC050000
0C000034
A88E0001
E1C27000
D4022004
A8630001
D4147008
D40E1804
040002F0
A8720000
03FFFF29
9D620008
0C000091
9CC5005B
BC450054
10000105
BC450154
B8AE004C
9CC5006E
03FFFF41
E0A63000
BC440004
0C00008B
BC440014
10000118
BC440054
9CC4005B
E0E63000
19600000
B8E70002
A96B9254
E0E75800
84870008
E4243800
0C0000FB
B8C60082
84C40004
9D60FFFC
E0C65803
E4833000
0C000006
15000000
84840008
E4272000
13FFFFF8
15000000
84E4000C
84740004
D402380C
D4022008
D4071008
03FFFF65
D404100C
1BC00000
18800000
ABDE924C
A8849ADC
847E0000
86C40000
BC23FFFF
0C0000EE
E2CEB000
9ED6100F
9CC0F000
E2D63003
A8720000
04000A69
A8960000
BC2BFFFF
0C000014
AB4B0000
19600000
E062C000
A96B9254
E443D000
E0825805
E0A02002
E0852004
9CA00001
B884005F
0C000079
D4012000
A4A500FF
BC050000
10000077
84810000
BC240000
0C000075
1B800000
84540008
9CE0FFFC
84A20004
E0A53803
E0657002
BDA3000F
10000003
9C800001
9C800000
A48400FF
BC240000
10000009
E44E2800
10000003
9CA00001
A8A40000
A4A500FF
BC050000
13FFFF98
A88E0001
0400028B
A8720000
03FFFEC4
9D600000
A86E0001
E1C27000
D4021804
A8A40001
D4147014
D4147010
E06E2000
D40E400C
D40E4008
D40E2804
D4032000
0400027C
A8720000
03FFFEB5
9D620008
03FFFF18
84740004
9C620008
84420014
E4031000
13FFFEEF
9CA50002
03FFFE9F
84820004
A8CE0001
8462000C
84A20008
D4023004
D405180C
E1C27000
03FFFFE5
D4032808
E0821800
84C2000C
84A40004
84E20008
A8A50001
A8720000
D4042804
D407300C
0400025F
D4063808
03FFFE98
9D620008
03FFFEB7
E0A63000
03FFFF60
A8A40000
B8830046
9CC40038
03FFFF79
E0E63000
856B0000
E40B1000
0C0000B6
15000000
A4650003
9C4BFFF8
BC230000
13FFFFF9
9CA5FFFF
84540004
AC66FFFF
E0431003
D4141004
E0C63000
E4A61000
10000003
9C600001
9C600000
A46300FF
BC030000
13FFFF37
E0603002
E0633004
BD630000
13FFFF33
E0623003
BC230000
13FFFEED
A8AD0000
E0C63000
E0623003
BC030000
13FFFFFD
9CA50004
03FFFEE7
E1652800
03FFFF89
9CA00000
1B800000
E423D000
AB9C9AAC
849C0000
E0962000
0C000066
D41C2000
84BE0000
BC25FFFF
0C000070
E07A1802
E0841800
D41C2000
A47A0007
BC030000
10000006
9CA01000
E35A1802
9CA01008
9F5A0008
E0A51802
E09AB000
A8720000
A4840FFF
E2C52002
040009C7
A8960000
BC0BFFFF
1000005B
9C600001
E06BD002
E0761800
A8630001
849C0000
84A10000
E0962000
D414D008
D41A1804
BC050000
10000011
D41C2000
BC58000F
0C000025
9CC0FFF8
84A20004
9C78FFF4
A4A50001
E0633003
9CE00005
E0A32804
E0C21800
D4022804
D4063804
BCA3000F
0C000047
D4063808
18400000
A8429AD8
84620000
E4A41800
10000003
18600000
D4022000
A8639AD4
84430000
E4441000
0C00001F
84540008
84A20004
9D60FFFC
D4032000
03FFFF4B
E0A55803
10000010
BC450554
B8AE004F
9CC50077
03FFFE3C
E0A63000
9C400001
03FFFF52
D41A1004
9CE00001
84740004
E0C73008
A8E40000
E0661804
03FFFF0E
D4141804
1000001B
15000000
B8AE0052
9CC5007C
03FFFE2C
E0A63000
03FFFF17
9ED60010
84A20004
9CE0FFFC
03FFFF2F
E0A53803
1000001F
BC440154
B883004C
9CC4006E
03FFFEE8
E0E63000
A4A30FFF
BC250000
13FFFF9A
15000000
E056C000
84740008
A8420001
03FFFFC6
D4031004
9CA000FC
03FFFE14
9CC0007E
03FFFFAA
9EC00000
18600000
A863924C
03FFFF92
D403D000
9C820008
18400000
A8720000
040005C1
A8429AAC
03FFFFB6
84820000
10000006
BC440554
B883004F
9CC40077
03FFFEC9
E0E63000
10000005
B8830052
9CC4007C
03FFFEC4
E0E63000
9CE000FC
03FFFEC1
9CC0007E
03FFFF55
84540004
A4C30003
D7E10FF8
D7E117FC
BC060000
9C21FFF8
1000004C
A4C400FF
BC050000
1000004B
9D65FFFF
8CA30000
E4053000
0C00000C
9C630001
9C63FFFF
00000026
9C210008
1000001F
15000000
8CA30000
E4253000
0C00001F
9D6BFFFF
9C630001
A4A30003
BC250000
13FFFFF7
BC0B0000
BCAB0003
0C00001C
BC0B0000
10000011
15000000
8C830000
E4043000
10000011
9C830001
00000006
E1635800
8CA4FFFF
E4253000
0C00000B
15000000
E4245800
A8640000
13FFFFFA
9C840001
9D600000
9C210008
8421FFF8
44004800
8441FFFC
9C210008
A9630000
8421FFF8
44004800
8441FFFC
A48400FF
B8A40008
E0852004
B8A40010
E0A52004
84830000
1840FEFE
E0852005
A842FEFF
E0E41000
AC84FFFF
18408080
E0872003
A8428080
E0841003
BC240000
13FFFFD6
BC0B0000
9D6BFFFC
BC4B0003
13FFFFF1
9C630004
03FFFFD0
BC0B0000
03FFFFCB
A9650000
03FFFFDD
A9650000
D7E10FF8
D7E117FC
BCA5000F
1000004C
9C21FFF8
E0C32004
A4C60003
BC260000
1000003B
A8C30000
9EE5FFF0
9CC40004
BAF70044
9E630004
9E240008
B9770004
9DE30008
9DA4000C
9D6B0014
9D83000C
E1645800
A9040000
A8E30000
86A80000
9CC60010
D407A800
E4265800
86A6FFF0
9D080010
D413A800
9CE70010
86B10000
9E730010
D40FA800
9E310010
86AD0000
9DEF0010
D40CA800
9DAD0010
13FFFFF0
9D8C0010
9CF70001
A565000F
B8E70004
BCAB0003
E0C33800
10000027
E0843800
A9860000
A9040000
A8EB0000
85A80000
9CE7FFFC
D40C6800
BC470003
9D8C0004
13FFFFFB
9D080004
9CEBFFFC
9C40FFFC
A4A50003
E0E71003
BC250000
9CE70004
E0C63800
0C000009
E0843800
E0A62800
8C440000
9CC60001
DBE617FF
E4262800
13FFFFFC
9C840001
9C210008
A9630000
8421FFF8
44004800
8441FFFC
A8C30000
BC250000
13FFFFF2
15000000
03FFFFF8
9C210008
03FFFFFB
A8AB0000
D7E10FF8
D7E117FC
E4A32000
10000015
9C21FFF8
E0C42800
E4633000
10000012
BCA5000F
E0832800
BC250000
0C000008
E0A42802
9CC6FFFF
8C460000
9C84FFFF
E4242800
13FFFFFC
D8041000
9C210008
A9630000
8421FFF8
44004800
8441FFFC
BCA5000F
0C000012
E0C32004
A8C30000
BC050000
13FFFFF6
15000000
E0A62800
8C440000
9CC60001
DBE617FF
E4262800
13FFFFFC
9C840001
9C210008
A9630000
8421FFF8
44004800
8441FFFC
A4C60003
BC260000
13FFFFF2
A8C30000
9EE5FFF0
9CC40004
BAF70044
9E630004
9E240008
BAB70004
9DE30008
9DA4000C
9EB50014
9D83000C
E2A4A800
A9040000
A8E30000
85680000
9CC60010
D4075800
E426A800
8566FFF0
9D080010
D4135800
9CE70010
85710000
9E730010
D40F5800
9E310010
856D0000
9DEF0010
D40C5800
9DAD0010
13FFFFF0
9D8C0010
9CF70001
A5A5000F
B8E70004
BCAD0003
E0C33800
10000014
E0843800
A9860000
A9040000
A8ED0000
85680000
9CE7FFFC
D40C5800
BC470003
9D8C0004
13FFFFFB
9D080004
9CEDFFFC
9C40FFFC
A4A50003
E0E71003
9CE70004
E0C63800
03FFFFB7
E0843800
03FFFFB5
A8AD0000
A4C30003
D7E10FF8
D7E117FC
BC060000
10000054
9C21FFF8
BC250000
0C00004C
9CA5FFFF
B9A40018
A8E30000
A8C30000
00000005
B9AD0098
BC050000
10000044
A8AC0000
9CC60001
D8076800
A5060003
9D85FFFF
BC280000
13FFFFF8
9CE70001
BCA50003
10000030
BC050000
A4E400FF
BCA5000F
B9070008
E0E83804
B9070010
1000001B
E0E83804
9E25FFF0
9D060004
BA310044
9DE60008
9DA6000C
B9710004
A9860000
9D6B0014
E1665800
D40C3800
D4083800
9D080010
D40F3800
D40D3800
E4285800
9D8C0010
9DEF0010
13FFFFF8
9DAD0010
9E310001
A4A5000F
BA310004
BCA50003
1000000F
E0C68800
A9860000
A9050000
9D08FFFC
D40C3800
BC480003
13FFFFFD
9D8C0004
9CE5FFFC
9C40FFFC
A4A50003
E0E71003
9CE70004
E0C63800
BC050000
1000000A
15000000
B8840018
E0A62800
B8840098
D8062000
9CC60001
E4262800
13FFFFFD
15000000
9C210008
A9630000
8421FFF8
44004800
8441FFFC
03FFFFC0
A8C30000
D7E117F0
18400000
D7E177F4
D7E197F8
D7E14FFC
D7E10FEC
9C21FFEC
A8429AE8
04000881
A9C30000
84620000
E4237000
0C00000C
AA4B0000
84820000
BC240000
13FFFFFE
18600000
A8AE0000
0400089D
A8639AE8
BC2B0000
13FFFFF8
15000000
18400000
A8429AE4
84620000
BC030000
0C000004
18600000
A8639AEC
D4039000
84620000
9C630001
D4021800
9C210014
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
18600000
D7E14FFC
A8639AE4
D7E10FF8
84830000
9C21FFF8
9C84FFFF
D4032000
84830000
BC240000
10000009
18600000
18A00000
A8639AEC
A8A59AE8
84630000
D4052000
0400085C
15000000
9C210008
8521FFFC
44004800
8421FFF8
D7E197E0
D7E1A7E4
D7E1C7EC
D7E14FFC
D7E10FD4
D7E117D8
D7E177DC
D7E1B7E8
D7E1D7F0
D7E1E7F4
D7E1F7F8
BC240000
9C21FFD4
AA440000
AB030000
0C0000B1
AA850000
07FFFFAE
9C54000B
84D2FFFC
9C60FFFC
BCA20016
9ED2FFF8
0C000052
E1C61803
9C800010
9CA00000
A8440000
E482A000
10000003
9C600001
9C600000
A46300FF
BC230000
100000A9
BC050000
0C0000A7
E56E2000
10000048
1B800000
E0767000
AB9C9254
84BC0008
E4051800
100000B5
9CE0FFFE
87830004
E0BC3803
E0A32800
84A50004
A4A50001
BC050000
0C000055
9CA0FFFC
E39C2803
E0BC7000
E5652000
1000008B
15000000
A4C60001
BC060000
0C000063
9CE0FFFC
8752FFF8
E356D002
84DA0004
E0C63803
E3853000
E57C2000
1000008A
9CAEFFFC
E3867000
E59C2000
10000058
A8940000
847A000C
849A0008
9CAEFFFC
D404180C
D4032008
BC450024
10000089
9C7A0008
BCA50013
1000000A
A8830000
84920000
BC45001B
D41A2008
84920004
100000E8
D41A200C
9C9A0010
9E520008
84B20000
AA830000
D4042800
A9DC0000
84720004
AADA0000
D4041804
84720008
D4041808
00000008
84DA0004
9C80FFF8
E0422003
A8820000
03FFFFB0
B8A2005F
AA920000
E06E1002
BCA3000F
0C000021
A4C60001
E0767000
E1C67004
D4167004
84430004
A8420001
D4031004
07FFFF70
A8780000
A9740000
9C21002C
8521FFFC
8421FFD4
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
A4C60001
BC060000
0C000015
9C60FFFC
8752FFF8
E356D002
84DA0004
03FFFFB7
E0C61803
E0961000
E0461004
A8A30001
D4161004
D4042804
E0441800
A8780000
84A20004
9C840008
A8A50001
04000361
D4022804
03FFFFDB
15000000
A8940000
07FFFB4D
A8780000
BC2B0000
0FFFFFD5
AA8B0000
84D2FFFC
9CA0FFFE
9C8BFFF8
E0662803
E0761800
E4241800
0C000090
9CAEFFFC
BC450024
1000007F
BCA50013
0C000068
BC45001B
A84B0000
A8720000
84830000
D4022000
84830004
D4022004
84630008
D4021808
A8920000
04000341
A8780000
03FFFFBB
15000000
07FFFB2E
A8850000
03FFFFBB
9C21002C
8483000C
84630008
AA920000
D403200C
D4041808
03FFFFA6
A9C50000
9C40000C
9D600000
03FFFFAF
D4181000
8483000C
84630008
D403200C
D4041808
847A000C
849A0008
BC450024
D404180C
D4032008
0FFFFF7B
9C7A0008
A8920000
07FFFE21
AA830000
A9DC0000
84DA0004
03FFFF90
AADA0000
87C50004
9CE0FFFC
9C620010
E3DE3803
E3DE7000
E57E1800
1000003A
A4C60001
BC060000
0FFFFFB6
9CA0FFFC
8752FFF8
E356D002
84DA0004
E0C62803
E3DE3000
E5A3F000
0FFFFF55
9CAEFFFC
847A000C
849A0008
D404180C
D4032008
BC450024
10000060
9E9A0008
BCA50013
1000000A
A8740000
84720000
BC45001B
D41A1808
84720004
1000005C
D41A180C
9C7A0010
9E520008
84920000
D4032000
84920004
D4032004
84920008
D4032008
E07E1002
E09A1000
A8630001
D41C2008
D4041804
A8780000
849A0004
A4840001
E0422004
07FFFED4
D41A1004
03FFFF65
A9740000
84520000
D40B1000
84520004
10000017
D40B1004
9C4B0008
03FFFF96
9C720008
E3DE1002
E2D61000
A87E0001
D41CB008
D4161804
A8780000
8492FFFC
A4840001
E0422004
07FFFEBF
D7F217FC
03FFFF50
A9720000
A86B0000
07FFFDCD
A8920000
03FFFF8B
A8920000
84520008
BC050024
D40B1008
8452000C
10000014
D40B100C
9C4B0010
03FFFF7B
9C720010
846BFFFC
9CE0FFFC
AA920000
E0633803
03FFFF2F
E1CE1800
84920008
BC050024
D41A2010
8492000C
1000000C
D41A2014
9C9A0018
03FFFF15
9E520010
84720010
9C4B0018
D40B1810
9C720018
84920014
03FFFF65
D40B2014
84B20010
9C9A0020
D41A2818
9E520018
84B2FFFC
03FFFF07
D41A281C
A8740000
07FFFDA2
A8920000
03FFFFB1
E07E1002
84720008
BC050024
D41A1810
8472000C
10000005
D41A1814
9C7A0018
03FFFFA1
9E520010
84920010
9C7A0020
D41A2018
9E520018
8492FFFC
03FFFF9A
D41A201C
D7E117F8
A8440000
9884000E
D7E14FFC
D7E10FF4
0400045B
9C21FFF4
BD8B0000
1000000A
9C80EFFF
84620050
E0635800
D4021850
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
9462000C
E0632003
DC02180C
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E10FFC
9C21FFFC
9D600000
9C210004
44004800
8421FFFC
98E4000C
D7E117EC
A8440000
A4870100
D7E177F0
D7E197F4
D7E1A7F8
D7E14FFC
D7E10FE8
BC040000
9C21FFE8
AA830000
AA450000
10000007
A9C60000
9882000E
9CA00000
0400041C
9CC00002
98E2000C
9C60EFFF
9882000E
E0E71803
A8B20000
DC02380C
A8740000
0400039C
A8CE0000
9C210018
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
D7E117F8
A8440000
9884000E
D7E14FFC
D7E10FF4
04000404
9C21FFF4
BC2BFFFF
0C00000A
9462000C
A8631000
D4025850
DC02180C
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
9C80EFFF
E0632003
DC02180C
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
9884000E
D7E14FFC
D7E10FF8
040003A1
9C21FFF8
9C210008
8521FFFC
44004800
8421FFF8
D7E117F4
D7E177F8
D7E14FFC
D7E10FF0
9C21FFF0
A9C30000
07FFFA11
A8440000
BC0B0000
10000006
15000000
846B0038
BC230000
0C000044
15000000
98A2000C
A485FFFF
A4640008
BC030000
10000018
A4640010
84C20010
BC260000
0C000021
A4640280
A4640001
BC030000
10000026
A4840002
84620014
9C800000
E0601802
D4022008
D4021818
BC260000
0C000026
9D600000
9C210010
8521FFFC
8421FFF0
8441FFF4
44004800
85C1FFF8
BC230000
0C00003C
A4840004
BC240000
10000026
15000000
84C20010
A8850008
BC260000
DC02200C
13FFFFE4
A484FFFF
A4640280
BC030200
13FFFFE1
A4640001
A8820000
040002BC
A86E0000
9482000C
03FFFFDA
84C20010
BC240000
10000003
15000000
84620014
D4021808
BC260000
13FFFFDE
9D600000
9862000C
A4830080
E4045800
13FFFFD9
A8630040
9D60FFFF
03FFFFD6
DC02180C
07FFF7B2
A86B0000
03FFFFBD
98A2000C
84820030
BC040000
1000000A
9C620040
E4041800
10000006
9C600000
040001CC
A86E0000
98A2000C
9C600000
D4021830
84C20010
9C80FFDB
9C600000
E0A52003
D4021804
03FFFFCC
D4023000
9C600009
A8A50040
D40E1800
DC02280C
03FFFFB9
9D60FFFF
D7E177F4
D7E14FFC
D7E10FEC
D7E117F0
D7E197F8
BC240000
9C21FFEC
0C00000D
A9C30000
BC030000
10000006
A8440000
84830038
BC240000
0C00003F
15000000
9862000C
BC030000
0C00000A
A86E0000
9C210014
9D600000
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
04000049
A8820000
AA4B0000
8562002C
BC0B0000
10000007
A86E0000
48005800
8482001C
BD6B0000
0C00002B
15000000
9462000C
A4630080
BC030000
0C000028
A86E0000
84820030
BC040000
10000009
9C620040
E4041800
10000005
9C600000
04000186
A86E0000
9C600000
D4021830
84820044
BC040000
10000006
15000000
0400017E
A86E0000
9C600000
D4021844
07FFF761
15000000
9C600000
07FFF763
DC02180C
9C210014
A9720000
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
07FFF748
15000000
03FFFFC2
9862000C
03FFFFD7
9E40FFFF
04000167
84820010
03FFFFD9
84820030
D7E14FFC
D7E117F8
D7E10FF4
9C21FFF4
07FFF94E
A8430000
A8820000
07FFFFA2
A86B0000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E117EC
9844000C
D7E1A7F8
AA830000
A462FFFF
D7E177F0
A9C40000
A4830008
D7E14FFC
D7E10FE8
D7E197F4
BC240000
10000044
9C21FFE8
A8420800
846E0004
BD430000
0C0000A3
DC0E100C
856E0028
BC0B0000
10000073
A442FFFF
9C600000
A4A21000
86540000
A4A5FFFF
E4051800
1000009E
D4141800
84AE0050
A4420004
BC020000
1000000A
A8740000
846E0030
844E0004
BC030000
10000004
E0A51002
844E003C
E0A51002
A8740000
848E001C
48005800
9CC00000
BC2BFFFF
0C000062
9C60F7FF
984E000C
848E0010
E0421803
D40E2000
A4621000
DC0E100C
9C400000
E4231000
10000079
D40E1004
848E0030
BC040000
1000004B
D4149000
9C4E0040
E4041000
10000004
15000000
04000112
A8740000
9C800000
D40E2030
9C210018
A9640000
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
864E0010
BC120000
10000036
A4630003
844E0000
BC230000
D40E9000
E0429002
10000003
9C600000
846E0014
BDA20000
0C000007
D40E1808
0000002B
9D600000
BD420000
0C000028
9D600000
A8B20000
A8C20000
856E0024
A8740000
48005800
848E001C
BD4B0000
E0425802
13FFFFF5
E2525800
944E000C
A8420040
9D60FFFF
DC0E100C
9C210018
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
84540000
BC220000
0C000046
AC620016
E0801802
E0641804
BD630000
10000007
AC42001D
E0601002
E0431004
BD820000
13FFFFE8
15000000
D4149000
9D600000
9C210018
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
84940000
AC44001D
E0602002
E0A01002
E0632004
E0451004
AC63FFFF
AC42FFFF
B863005F
B842005F
E0431004
BC220000
10000007
AC840016
E0402002
E0822004
BD640000
0C000022
15000000
984E000C
9C80F7FF
84AE0010
E0422003
D40E2800
A4821000
DC0E100C
9C400000
E4241000
0FFFFF8E
D40E1004
BC230000
0FFFFF8B
15000000
03FFFF89
D40E5850
846E003C
BD430000
13FFFF5D
9D600000
03FFFFD2
9C210018
A8740000
848E001C
48005800
9CC00001
BC2BFFFF
0FFFFFBA
A8AB0000
944E000C
03FFFF5D
856E0028
944E000C
A8420040
03FFFFAB
DC0E100C
D7E117F4
D7E177F8
D7E14FFC
D7E10FF0
BC030000
9C21FFF0
A8430000
10000006
A9C40000
84830038
BC240000
0C00000F
15000000
986E000C
BC030000
10000005
9D600000
A8620000
07FFFF26
A88E0000
9C210010
8521FFFC
8421FFF0
8441FFF4
44004800
85C1FFF8
07FFF64E
15000000
03FFFFF2
986E000C
D7E117F8
D7E14FFC
D7E10FF4
BC230000
9C21FFF4
0C00000C
A8430000
07FFF857
15000000
A8820000
07FFFFD8
A86B0000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
18400000
18800000
A8426DF4
A88453E8
07FFF814
84620000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E1A7F8
1A800000
D7E117EC
D7E177F0
D7E197F4
D7E14FFC
D7E10FE8
9C21FFE8
AA949254
A8440000
07FFFC0B
AA430000
84740008
85C30004
9C60FFFC
E1CE1803
9C60F000
E04E1002
9C420FEF
E0421803
E0421800
BD420FFF
0C000009
A8720000
040003DA
9C800000
84740008
E0637000
E42B1800
0C00000D
A8720000
07FFFC20
A8720000
9C210018
9D600000
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
040003C8
E0801002
BC2BFFFF
0C000015
18800000
E1CE1002
A8849AAC
84B40008
84640000
A9CE0001
E0431002
D4057004
A8720000
07FFFC08
D4041000
9C210018
9D600001
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
A8720000
040003AF
9C800000
84740008
E04B1802
BDA2000F
13FFFFD7
18800000
A8420001
A884924C
D4031004
84840000
18400000
E16B2002
A8429AAC
03FFFFCE
D4025800
D7E177F8
D7E14FFC
D7E10FF0
D7E117F4
BC040000
9C21FFF0
1000004F
A9C30000
07FFFBBA
A8440000
8462FFFC
9C80FFFE
19000000
E0A32003
9CE2FFF8
A9089254
E0C72800
85680008
84860004
E42B3000
9D60FFFC
A4630001
0C000063
E0845803
BC230000
1000000E
D4062004
8442FFF8
18600000
E0E71002
E0A51000
A863925C
84470008
E4021800
10000070
15000000
8467000C
D402180C
D4031008
E0462000
84420004
A4420001
BC020000
0C000011
A8650001
E0A52000
18800000
84460008
A884925C
E4022000
10000081
A8850001
8486000C
A8650001
D402200C
D4041008
E0472800
D4071804
00000005
D4022800
E0472800
D4071804
D4022800
BC4501FF
1000001B
B8450049
B8A50043
9C800001
84680004
E0452800
B8A50082
B8420002
E0A42808
18800000
A8849254
E0A51804
E0422000
D4082804
84820008
D407100C
D4072008
D4023808
D404380C
07FFFB99
A86E0000
9C210010
8521FFFC
8421FFF0
8441FFF4
44004800
85C1FFF8
BC420004
1000004A
BC420014
B8450046
9C620038
E0431800
19600000
B8420002
A96B9254
E0425800
84820008
E4241000
0C000044
15000000
84C40004
9C60FFFC
E0C61803
E4462800
0C000006
15000000
84840008
E4222000
13FFFFF8
15000000
84A4000C
D407280C
D4072008
D4053808
03FFFFDC
D404380C
BC230000
10000009
E0A42800
8442FFF8
E0E71002
E0A51000
84670008
8447000C
D403100C
D4021808
18400000
A8650001
A8429250
D4071804
84420000
E4651000
0FFFFFCA
D4083808
18400000
A86E0000
A8429ADC
07FFFF1F
84820000
03FFFFC3
15000000
E0462000
84420004
A4420001
BC020000
0C00000C
E0472800
8446000C
84660008
E0852000
D403100C
A8A40001
D4021808
E0472000
D4072804
03FFFFB3
D4022000
A8650001
D4071804
03FFFFAF
D4022800
10000015
BC420054
9C62005B
03FFFFB8
E0431800
B8430082
9C600001
84C80004
E0431008
A8A40000
E0423004
03FFFFC3
D4081004
D4083814
D4083810
E0672800
D407100C
D4071008
D4072004
03FFFF9A
D4032800
10000006
BC420154
B845004C
9C62006E
03FFFFA2
E0431800
10000006
BC420554
B845004F
9C620077
03FFFF9C
E0431800
10000006
15000000
B8450052
9C62007C
03FFFF96
E0431800
9C4000FC
03FFFF93
9C60007E
98A4000C
A4C5FFFF
D7E117EC
A4460002
D7E177F0
D7E14FFC
D7E10FE8
D7E197F4
D7E1A7F8
BC020000
9C21FFAC
0C00003B
A9C30000
A8440000
9884000E
BD840000
10000018
A4C60080
040000AC
A8A10000
BD6B0000
0C000010
84810004
A8A08000
A484F000
AC642000
E4242800
E2401802
E2521804
AE52FFFF
0C000037
BA52005F
9462000C
A8630800
9E800400
0000000B
DC02180C
98A2000C
A4C5FFFF
A4C60080
BC060000
0C00002A
9E800400
A8A50800
9E400000
DC02280C
A86E0000
07FFF6F2
A8940000
BC2B0000
0C000039
18800000
9462000C
A8630080
A88429C4
BC120000
D40E203C
DC02180C
D4025800
D4025810
0C000025
D402A014
9C210054
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
9C440043
D4041000
D4041010
9C400001
D4041014
9C210054
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
03FFFFD8
9E800040
18800000
84620028
A8844CF0
E4232000
13FFFFC7
15000000
9462000C
9E800400
E063A004
D402A04C
03FFFFCF
DC02180C
9882000E
04000074
A86E0000
BC0B0000
13FFFFD9
15000000
9462000C
A8630001
03FFFFD5
DC02180C
9862000C
A4830200
BC040000
0FFFFFD0
A8630002
9C820043
DC02180C
9C600001
D4022000
D4022010
03FFFFC9
D4021814
D7E117F0
D7E177F4
D7E197F8
D7E14FFC
D7E10FEC
BC260000
9C21FFEC
AA460000
A8450000
10000009
E1C53000
00000014
9C210014
0400010A
9C420001
E4227000
0C00000E
15000000
90620000
BC23000A
13FFFFF9
15000000
9C60000D
04000100
9C420001
040000FE
9062FFFF
E4227000
13FFFFF6
15000000
9C210014
A9720000
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
D7E14FFC
D7E10FF8
040003F9
9C21FFF8
15000000
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E14FFC
D7E10FF8
040003EA
9C21FFF8
9C600058
D40B1800
9C210008
9D60FFFF
8521FFFC
44004800
8421FFF8
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800058
9C210004
9D600000
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E14FFC
D7E10FF8
040003AF
9C21FFF8
9C600058
D40B1800
9C210008
9D60FFFF
8521FFFC
44004800
8421FFF8
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800005
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800005
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
18600000
D7E10FFC
A8636BB0
9C21FFFC
84630000
9C630002
8C630000
9C210004
44004800
8421FFFC
D7E117F4
18400000
D7E177F8
A8426BB0
D7E14FFC
85C20000
D7E10FF0
BC0E0000
1000002C
9C21FFF0
18600000
18A00000
A8636BB4
9CC00000
84830000
18600000
A8A59AF0
A8636BAC
B8840004
84630000
D4053000
04000367
9DCE0003
9C60FF80
A48B00FF
D80E1800
A56BFFFF
84620000
9CC0FFC3
D8032000
B86B0048
84820000
9D600000
9C840001
D8041800
9C800003
84620000
9C630003
D8032000
84620000
9C630002
D8033000
9C600000
84420000
9C420001
D8021800
9C210010
8521FFFC
8421FFF0
8441FFF4
44004800
85C1FFF8
03FFFFFA
9D60FFFF
18800000
B8630018
A8846BB0
D7E10FFC
84C40000
B8630098
9C21FFFC
9CA60005
8C850000
A4840020
BC040000
13FFFFFD
15000000
A46300FF
D8061800
9C210004
44004800
8421FFFC
D7E117F8
18400000
D7E14FFC
A8426BB0
D7E10FF4
84820000
18400000
9C840001
A8429AF0
9C21FFF4
D4021800
9C400001
9CA00000
D8041000
18400000
18800000
A8426BB8
A8845DE0
040000DF
84620000
04000133
84620000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
18800000
A8846BB0
84840000
E4040000
10000004
15000000
03FFFFCD
15000000
44004800
15000004
B4600001
A4830004
E4040000
10000021
15000000
B4C00011
9CA0FFFF
ACA50010
E0A62803
C0002811
B4600006
A4830080
B8E40047
A9000010
E1C83808
A4830078
B8E40043
A9000001
E1A83808
9CC00000
E0AE3808
C0803002
E4262800
13FFFFFE
E0C67000
B4C00011
A8C60010
C0003011
15000000
15000000
15000000
15000000
15000000
15000000
15000000
15000000
B4600001
A4830002
E4040000
10000019
15000000
B4C00011
9CA0FFFF
ACA50008
E0A62803
C0002811
B4600005
A4830080
B8E40047
A9000010
E1C83808
A4830078
B8E40043
A9000001
E1A83808
9CC00000
E0AE3808
C0603003
E4262800
13FFFFFE
E0C67000
B4C00011
A8C60008
C0003011
44004800
15000000
B5A00011
A9AD0010
C0006811
15000000
15000000
15000000
15000000
15000000
44004800
15000000
B5A00011
9D80FFFF
AD8C0010
E18D6003
C0006011
44004800
15000000
44004800
C0801802
B5A00011
A9AD0008
C0006811
15000000
15000000
15000000
15000000
15000000
44004800
15000000
B5A00011
9D80FFFF
AD8C0008
E18D6003
C0006011
44004800
15000000
44004800
C0601803
D4011008
D4012814
D4013018
D401381C
D4014020
D4014824
D4015028
D401582C
D4016030
D4016834
D4017038
D401783C
D4018040
D4018844
D4019048
D401984C
D401A050
D401A854
D401B058
D401B85C
D401C060
D401C864
D401D068
D401D86C
D401E070
D401E874
D401F078
D401F87C
B5C00020
D4017080
B5C00040
D4017084
1A800000
AA949664
86940000
1AA00000
AAB59C04
D415A000
A5A3FF00
B9AD0046
9DADFFF8
19C00000
A9CE9C20
E1CE6800
85AE0000
E42D0000
0C000034
15000000
48006800
E0642004
1A800000
AA949C08
86940000
1AA00000
AAB59C04
D415A000
18400000
A8429C0C
84620000
9C63FFFF
D4021800
84410080
C0001020
84410084
C0001040
84410008
8461000C
84810010
84A10014
84C10018
84E1001C
85010020
85210024
85410028
8561002C
85810030
85A10034
85C10038
85E1003C
86010040
86210044
86410048
8661004C
86810050
86A10054
86C10058
86E1005C
87010060
87210064
87410068
8761006C
87810070
87A10074
87C10078
87E1007C
84210004
24000000
15000000
07FFF04A
E0642004
D7E117FC
18400000
B8630002
A8429AF4
D7E10FF8
E0C31000
18400000
9C21FFF8
A8429B74
D4062000
E0631000
D4032800
9C210008
8421FFF8
44004800
8441FFFC
D7E10FFC
9C800011
9C21FFFC
B4640000
A8630004
C0041800
9C210004
44004800
8421FFFC
D7E10FF8
D7E117FC
9C600011
9C21FFF8
B5630000
9C40FFFB
E08B1003
C0032000
9C210008
B96B0042
8421FFF8
A56B0001
44004800
8441FFFC
D7E10FF8
D7E117FC
9C800011
9C21FFF8
B4840000
9C40FFFB
BC230000
E0841003
10000003
9CA00004
A8A30000
E0652004
9C800011
C0041800
9C210008
8421FFF8
44004800
8441FFFC
9C21FFFC
D4014800
B6804802
1A000000
AA109AF4
1A400000
AA529B74
E094000F
E4240000
0C000010
15000000
9EC4FFFF
B8D60002
E1C68000
E1A69000
85CE0000
E42E0000
0C000004
15000000
48007000
846D0000
A8C00001
E0C6B008
03FFFFF0
E2943005
85210000
C120A002
44004800
9C210004
9C21FFFC
D4012000
A8800001
E0841808
B4604800
E0632004
C1201800
84810000
44004800
9C210004
9C21FFFC
D4012000
A8800001
E0841808
AC84FFFF
B4604800
E0632003
C1201800
84810000
44004800
9C210004
D7E14FFC
D7E117E4
D7E197EC
D7E1A7F0
D7E1B7F4
D7E1C7F8
D7E10FE0
D7E177E8
9C21FFE0
AA840000
07FFFFA4
18400000
04000170
AACB0000
18600000
A8429660
A8639BF4
9C800000
84A20000
AB0B0000
040000BF
AA430000
84520000
18600000
A8820000
A8639BF4
040000B9
E0B41000
E42B1000
13FFFFF9
A9CB0000
0400016B
A8780000
07FFFF9B
A8760000
9C210020
A96E0000
8521FFFC
8421FFE0
8441FFE4
85C1FFE8
8641FFEC
8681FFF0
86C1FFF4
44004800
8701FFF8
D7E117D8
18400000
D7E1F7F8
A8428E24
9FC00424
D7E14FFC
D7E177DC
D7E197E0
D7E1A7E4
D7E1B7E8
D7E1C7EC
D7E1D7F0
D7E1E7F4
84620000
A8BE0000
D7E10FD4
9C800000
9C21FFD4
07FFF789
1B400000
84C20000
1B800000
9C860354
9C6603BC
9CA602EC
AB5A6DF8
9F00330E
9EC0ABCD
9E801234
9E40E66D
9DC0DEEC
AB9C9664
D4062008
D406180C
9C80000B
9C600005
D4062804
D406D034
DC06C0AC
DC06B0AE
DC06A0B0
DC0690B2
DC0670B4
DC0618B6
DC0620B8
847C0000
A8BE0000
9CE00000
9D000001
D40638A4
D40640A8
07FFF768
9C800000
847C0000
84420000
9C8303BC
9D000005
D403200C
9C80000B
DC0340B6
DC0320B8
18800000
9CC302EC
A8849C08
9CA30354
D4041000
18800000
9CE00000
A8849C04
9D000001
DC03C0AC
DC03B0AE
DC03A0B0
DC0390B2
DC0370B4
D40338A4
D40340A8
D403D034
D4041000
D4033004
D4032808
9C21002C
8521FFFC
8421FFD4
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
18600000
D7E10FFC
A8639C04
9C21FFFC
85630000
9C210004
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C210004
44004800
8421FFFC
D7E14FFC
D7E117F8
D7E10FF4
9C21FFF4
07FFFFF7
9C400000
18800000
18600000
A88463D0
A8639C20
D4032018
18600000
A8639C0C
D4031000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E14FFC
D7E117F8
D7E10FF4
07FFFEFF
9C21FFF4
040000CB
A84B0000
9C21000C
E0421000
8521FFFC
8421FFF4
E1625804
44004800
8441FFF8
D7E14FFC
D7E117F8
D7E10FF4
A8430000
9C21FFF4
040000CB
A4630001
B8620041
07FFFEFA
A4630001
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
44004800
E1600004
44004800
E1600004
44004800
A9600001
44004800
85630000
44004800
D4032000
85630000
E40B2000
0C000003
15000000
D4032800
44004800
15000000
E0800004
03FFFFF8
9CA00001
9C63FFFE
D7E117FC
18400000
B8630002
A8429C20
D7E10FF8
E0631000
9C21FFF8
D4032000
9C210008
8421FFF8
44004800
8441FFFC
18A00000
D7E10FF8
A8A59BF8
D7E117FC
84650000
9C21FFF8
9C630001
9C805000
D4051800
B4640000
18402FFF
A842FFFF
E0631003
18406000
E0631004
C0041800
9C210008
8421FFF8
44004800
8441FFFC
D7E197F8
D7E14FFC
D7E10FEC
D7E117F0
D7E177F4
9E400001
9C21FFEC
B4B20000
B8A5004A
E0A59003
BC050000
10000020
18400000
A8830000
A8426BAC
19C00000
84620000
040000C9
18400FFF
A842FFFF
A9CE9BF8
E16B1003
9C405000
D40E5804
C0025800
18800000
9C400000
9C600005
A8846840
D40E1000
07FFFFC1
15000000
9C605001
D40E9008
C0031000
A9620000
9C210014
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
03FFFFF9
9D60FFFF
A8830000
18600000
D7E117F8
A8636BAC
18400FFF
D7E14FFC
D7E10FF4
84630000
9C21FFF4
040000A4
A842FFFF
9C805000
E16B1003
B4640000
1840F000
E0631003
E0635804
C0041800
18600000
A8639BF8
D4035804
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E14FFC
D7E10FF8
A8830000
9C21FFF8
07FFFF94
9C600005
9C210008
8521FFFC
44004800
8421FFF8
18800000
D7E10FF8
A8849BF8
D7E117FC
9CA05000
9C21FFF8
D4041808
B4850000
B8C4005E
BC060000
10000007
B863001E
18403FFF
A842FFFF
E0841003
E0641804
C0051800
9C210008
8421FFF8
44004800
8441FFFC
D7E10FF8
D7E117FC
9CA05000
9C21FFF8
B4650000
18403FFF
A842FFFF
E0831003
18600000
18402000
A8639BF8
84630008
B863001E
E0631004
E0632004
C0051800
9C800011
B4640000
A8630002
C0041800
9C210008
8421FFF8
44004800
8441FFFC
D7E10FF8
D7E117FC
9C600011
9C21FFF8
B5630000
9C40FFFD
E08B1003
C0032000
9C210008
B96B0041
8421FFF8
A56B0001
44004800
8441FFFC
D7E10FFC
9C800011
9C21FFFC
B4640000
A8630002
C0041800
9C210004
44004800
8421FFFC
D7E10FF8
D7E117FC
9C805000
9C21FFF8
B4640000
18403FFF
A842FFFF
E0631003
C0041800
9C210008
8421FFF8
44004800
8441FFFC
D7E10FF8
D7E117FC
9C805000
9C21FFF8
B4640000
1840EFFF
A842FFFF
E0631003
C0041800
9C800000
9C605001
C0032000
9C210008
8421FFF8
44004800
8441FFFC
18600000
D7E10FFC
A8639BF8
9C21FFFC
85630000
9C210004
44004800
8421FFFC
18600000
D7E117FC
A8639BF8
9C400000
D7E10FF8
9C21FFF8
D4031000
9C210008
8421FFF8
44004800
8441FFFC
04000000
02FAF080
90000000
0001C200
00000002
1500000C
15000000
44004800
15000000
44004800
15000000
D7E14FFC
D7E10FF8
07FFF27E
9C21FFF8
9C210008
8521FFFC
44004800
8421FFF8
9C21FFFC
D4014800
9D600000
9D040000
9CA30000
E4285800
0C000036
9CE00000
E4482800
10000032
E4082800
1000002E
E48B4000
0C00000D
9DA00020
19208000
9CC0FFFF
E0654803
B8870001
9DE50000
B863005F
E1AD3000
E0E41804
E4874000
13FFFFF9
B8A50001
B8E70041
9DAD0001
9D200000
E4896800
0C00001E
9CAF0000
19E08000
9E200000
E0657803
B8870001
B863005F
E0E41804
E0C74002
E0667803
B863005F
9C800000
E4232000
10000003
B86B0001
9C800001
B8A50001
E4248800
0C000003
E1632004
9CE60000
9D290001
E4896800
13FFFFED
15000000
00000005
15000000
00000003
9D600001
9CE50000
85210000
44004800
9C210004
9C21FFF8
D4014800
D4017004
9CA30000
9DC00000
E5850000
0C000004
9C600000
9DC00001
E0A02802
E5840000
0C000004
15000000
9DCE0001
E0802002
07FFFFB2
9C650000
BC0E0001
0C000003
15000000
E1605802
85210000
85C10004
44004800
9C210008
D7E117F8
18400000
D7E14FFC
A8428E08
D7E10FF4
8462FFFC
9C21FFF4
BC23FFFF
0C000008
9C42FFFC
48001800
9C42FFFC
84620000
BC23FFFF
13FFFFFC
15000000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E14FFC
D7E10FF8
9C21FFF8
9C210008
8521FFFC
44004800
8421FFF8
9C21FFFC
D4014800
07FFED0E
15000000
85210000
44004800
9C210004
48656C6C
6F20576F
726C6421
00008E28
43000A00
7FFFFFFF
FFFFFFFF
FFFFFFFF
00002000
00002000
00008E28
00009114
0000917C
000091E4
00006DF8
00000001
330EABCD
1234E66D
DEEC0005
000B0000
FFFFFFFF
00020000
00009254
00009254
0000925C
0000925C
00009264
00009264
0000926C
0000926C
00009274
00009274
0000927C
0000927C
00009284
00009284
0000928C
0000928C
00009294
00009294
0000929C
0000929C
000092A4
000092A4
000092AC
000092AC
000092B4
000092B4
000092BC
000092BC
000092C4
000092C4
000092CC
000092CC
000092D4
000092D4
000092DC
000092DC
000092E4
000092E4
000092EC
000092EC
000092F4
000092F4
000092FC
000092FC
00009304
00009304
0000930C
0000930C
00009314
00009314
0000931C
0000931C
00009324
00009324
0000932C
0000932C
00009334
00009334
0000933C
0000933C
00009344
00009344
0000934C
0000934C
00009354
00009354
0000935C
0000935C
00009364
00009364
0000936C
0000936C
00009374
00009374
0000937C
0000937C
00009384
00009384
0000938C
0000938C
00009394
00009394
0000939C
0000939C
000093A4
000093A4
000093AC
000093AC
000093B4
000093B4
000093BC
000093BC
000093C4
000093C4
000093CC
000093CC
000093D4
000093D4
000093DC
000093DC
000093E4
000093E4
000093EC
000093EC
000093F4
000093F4
000093FC
000093FC
00009404
00009404
0000940C
0000940C
00009414
00009414
0000941C
0000941C
00009424
00009424
0000942C
0000942C
00009434
00009434
0000943C
0000943C
00009444
00009444
0000944C
0000944C
00009454
00009454
0000945C
0000945C
00009464
00009464
0000946C
0000946C
00009474
00009474
0000947C
0000947C
00009484
00009484
0000948C
0000948C
00009494
00009494
0000949C
0000949C
000094A4
000094A4
000094AC
000094AC
000094B4
000094B4
000094BC
000094BC
000094C4
000094C4
000094CC
000094CC
000094D4
000094D4
000094DC
000094DC
000094E4
000094E4
000094EC
000094EC
000094F4
000094F4
000094FC
000094FC
00009504
00009504
0000950C
0000950C
00009514
00009514
0000951C
0000951C
00009524
00009524
0000952C
0000952C
00009534
00009534
0000953C
0000953C
00009544
00009544
0000954C
0000954C
00009554
00009554
0000955C
0000955C
00009564
00009564
0000956C
0000956C
00009574
00009574
0000957C
0000957C
00009584
00009584
0000958C
0000958C
00009594
00009594
0000959C
0000959C
000095A4
000095A4
000095AC
000095AC
000095B4
000095B4
000095BC
000095BC
000095C4
000095C4
000095CC
000095CC
000095D4
000095D4
000095DC
000095DC
000095E4
000095E4
000095EC
000095EC
000095F4
000095F4
000095FC
000095FC
00009604
00009604
0000960C
0000960C
00009614
00009614
0000961C
0000961C
00009624
00009624
0000962C
0000962C
00009634
00009634
0000963C
0000963C
00009644
00009644
0000964C
0000964C
00009AE0
00009C98
00009668
00009954
000099BC
00009A24
00006DF8
00000001
330EABCD
1234E66D
DEEC0005
000B0000
	 
