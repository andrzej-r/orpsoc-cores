@00000000
18000000
18400000
A8421000
18800400
A8841000
18609500
A8630000
84A30200
B8A50044
18609600
A8630000
D4032804
18600001
A8630203
D4021800
18600405
A8630607
D4021804
18600809
A8630A0B
D4021808
18600C0D
A8630E0F
D402180C
18601011
A8631213
D4041800
18601415
A8631617
D4041804
18601819
A8631A1B
D4041808
18601C1D
A8631E1F
D404180C
84E20000
84E20004
84E20008
84E2000C
84E40000
84E40004
84E40008
84E4000C
15000001
	 
