@00000000
18000000
18400000
A8421000
18A0FFFF
A8A5FFFF
18C09100
A8C62000
DC062804
18600001
A8630203
D4021800
18600405
A8630607
D4021804
18600000
A8630008
D8021808
18600000
A8630009
D8021809
18600000
A8630A0B
DC02180A
18600000
A8630C0D
DC02180C
18600000
A863000E
D802180E
18600000
A863000F
D802180F
18601011
A8631213
D4021810
18601415
A8631617
D4021814
18601819
A8631A1B
D4021818
18601C1D
A8631E1F
D402181C
18600000
A8630000
8C820000
E4032000
0C00003D
18600000
A8630001
8C820001
E4032000
0C000038
18600000
A8630203
94820002
E4032000
0C000033
18600000
A8630405
94820004
E4032000
0C00002E
18600000
A8630006
8C820006
E4032000
0C000029
18600000
A8630007
8C820007
E4032000
0C000024
18600809
A8630A0B
84820008
E4032000
0C00001F
18600C0D
A8630E0F
8482000C
E4032000
0C00001A
18601011
A8631213
84820010
E4032000
0C000015
18601415
A8631617
84820014
E4032000
0C000010
18601819
A8631A1B
84820018
E4032000
0C00000B
18601C1D
A8631E1F
8482001C
E4032000
0C000006
18A0FFFF
A8A5FFFF
DC062800
03FFFFFD
15000000
18A0DEAD
A8A5DEAD
DC062800
03FFFFFD
15000000
	 
