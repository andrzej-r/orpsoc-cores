@00000000
18000000
18200000
18400000
18600000
18800000
18A00000
18C00000
18E00000
19000000
19200000
19400000
19600000
19800000
19A00000
19C00000
19E00000
1A000000
1A200000
1A400000
1A600000
1A800000
1AA00000
1AC00000
1AE00000
1B000000
1B200000
1B400000
1B600000
1B800000
1BA00000
1BC00000
1BE00000
A8200001
C0000811
C1400000
18800000
A8842030
44002000
15000000
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003E97
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003E57
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003E17
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003DD7
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003D97
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003D57
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003D17
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003CD7
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003C97
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003C57
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003C17
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003BD7
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003B97
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003B57
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003B17
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003AD7
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003A97
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003A57
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003A17
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
000039D7
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003997
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003957
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003917
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
000038D7
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003897
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003857
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003817
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
000037D7
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003797
B4800020
D4000804
18200001
A8215134
84210000
E4010000
0C000006
15000000
18200001
A8215138
00000004
84210000
84200004
9C21FF80
9C21FF78
D401180C
84600004
D4011804
D4012010
18600001
A8635134
84830000
9C840001
D4032000
B4600010
00003757
B4800020
15000000
15000000
9C21FFFC
D4014800
040000BC
15000000
04003E7C
15000000
85210000
44004800
9C210004
44004800
15000000
040036BB
15000000
040039BC
15000000
18600001
A8634FA8
18800001
A88451C0
D4030000
E4832000
13FFFFFE
9C630004
18200001
A8210704
84210000
18400001
A8420708
84420000
E0211000
18600001
A8635138
D4030800
18600001
A86342A8
84630000
E0811802
18A00001
A8A55140
D4052000
E0202004
E0410804
18600001
A863513C
D4030800
18600001
A86342A4
84630000
E0811802
18A00001
A8A55144
D4052000
04003862
15000000
040037F5
15000000
07FFFFC8
15000000
18600001
04000AD1
A8631A74
18800001
A8840710
84840000
E4240000
0C000004
E0600004
04003616
15000000
04003986
15000000
E0600004
E0800004
0400023B
E0A00004
04000ACD
9C6B0000
15000000
D7E117F8
18600001
18400001
A8634FAB
A8424FA8
D7E14FFC
E0631002
D7E10FF4
BCA30006
10000009
9C21FFF4
18800000
A8840000
BC040000
10000004
15000000
48002000
A8620000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E117F8
18600001
18400001
A8634FA8
A8424FA8
D7E14FFC
E0631002
D7E10FF4
B8630082
B883005F
E0841800
B8840081
BC040000
10000009
9C21FFF4
18A00000
A8A50000
BC050000
10000004
15000000
48002800
A8620000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E197F8
1A400001
D7E117F0
AA524FA8
D7E14FFC
8C520000
D7E10FEC
D7E177F4
BC220000
10000026
9C21FFEC
19C00001
18800001
A9CE429C
A8844298
18400001
E1CE2002
A8424FAC
B9CE0082
84620000
9DCEFFFF
E4837000
0C00000E
9C630001
18A00001
B8830002
A8A54298
D4021800
E0642800
84630000
48001800
15000000
84620000
E4837000
13FFFFF6
9C630001
07FFFFAA
18400000
A8420000
BC220000
0C000006
9C400001
18600001
07FFF753
A863428C
9C400001
D8121000
9C210014
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
D7E14FFC
D7E10FF8
9C21FFF8
9C210008
8521FFFC
44004800
8421FFF8
18600000
D7E14FFC
A8630000
D7E10FF8
BC030000
10000007
9C21FFF8
18600001
18800001
A863428C
07FFF737
A8844FB0
18600001
A86342A0
84830000
BC040000
0C000008
18800000
07FFFF96
15000000
9C210008
8521FFFC
44004800
8421FFF8
A8840000
BC040000
13FFFFF8
15000000
48002000
15000000
03FFFFF4
15000000
D7E14FFC
D7E10FF8
9C21FFF8
9C210008
8521FFFC
44004800
8421FFF8
D7E117FC
9C410000
9C21FFEC
D7E21FEC
18609100
A8634000
9C800001
DC032000
9C600000
D7E21FF8
00000017
15000000
8482FFEC
8462FFF8
E0641848
A463000F
D7E21FF4
18800001
A88442B0
8462FFF4
E0641800
8C630000
D7E21FF0
8462FFF8
18809100
A884403C
E0641802
8482FFF0
A484FFFF
DC032000
8462FFF8
9C630004
D7E21FF8
8462FFF8
BDA3001F
13FFFFE9
15000000
A8220000
8441FFFC
44004800
15000000
D7E117F8
9C410000
D7E14FFC
D7E177F4
9C21FFD8
D7E21FE8
D7E227E4
8462FFE8
D7E21FF0
00000016
15000000
8462FFF0
8482FFF0
D4032000
8462FFF0
A46300FF
BC230000
1000000B
15000000
8462FFF0
07FFFFC3
15000000
8462FFF0
D4011800
18600001
A8631A90
04000A0D
15000000
8462FFF0
9C630004
D7E21FF0
8482FFF0
8462FFE4
E4841800
13FFFFE9
15000000
8462FFE8
D7E21FF0
00000025
15000000
8462FFF0
84630000
D7E21FEC
8462FFF0
A46300FF
BC230000
1000000B
15000000
8462FFF0
07FFFFA6
15000000
8462FFF0
D4011800
18600001
A8631AA7
040009F0
15000000
8482FFEC
8462FFF0
E4041800
1000000C
15000000
8462FFEC
D4011800
8462FFF0
D4011804
8462FFF0
D4011808
18600001
A8631ABD
040009E1
15000000
8462FFF0
9C630004
D7E21FF0
8482FFF0
8462FFE4
E4841800
13FFFFDA
15000000
8462FFE8
D7E21FF0
0000001B
15000000
85C2FFF0
8462FFF0
A880FFFF
0400013C
15000000
A86B0000
A463FFFF
DC0E1800
8462FFF0
A46300FF
BC230000
1000000B
15000000
8462FFF0
07FFFF75
15000000
8462FFF0
D4011800
18600001
A8631AF2
040009BF
15000000
8462FFF0
9C630002
D7E21FF0
8482FFF0
8462FFE4
E4841800
13FFFFE4
15000000
8462FFE8
D7E21FF0
00000030
15000000
8462FFF0
94630000
A463FFFF
D7E21FEC
8462FFF0
A46300FF
BC230000
1000000B
15000000
8462FFF0
07FFFF57
15000000
8462FFF0
D4011800
18600001
A8631B09
040009A1
15000000
8462FFF0
A880FFFF
04000109
15000000
A86B0000
A8830000
8462FFEC
E4041800
10000011
15000000
8462FFF0
A880FFFF
040000FF
15000000
A86B0000
A8830000
8462FFEC
D4011800
8462FFF0
D4011804
D4012008
18600001
A8631B1F
04000988
15000000
8462FFF0
9C630002
D7E21FF0
8482FFF0
8462FFE4
E4841800
13FFFFCF
15000000
8462FFE8
D7E21FF0
0000001B
15000000
85C2FFF0
8462FFF0
9C8000FF
040000E3
15000000
A86B0000
A46300FF
D80E1800
8462FFF0
A46300FF
BC230000
1000000B
15000000
8462FFF0
07FFFF1C
15000000
8462FFF0
D4011800
18600001
A8631B54
04000966
15000000
8462FFF0
9C630001
D7E21FF0
8482FFF0
8462FFE4
E4841800
13FFFFE4
15000000
8462FFE8
D7E21FF0
00000030
15000000
8462FFF0
8C630000
A46300FF
D7E21FEC
8462FFF0
A46300FF
BC230000
1000000B
15000000
8462FFF0
07FFFEFE
15000000
8462FFF0
D4011800
18600001
A8631B6A
04000948
15000000
8462FFF0
9C8000FF
040000B0
15000000
A86B0000
A8830000
8462FFEC
E4041800
10000011
15000000
8462FFF0
9C8000FF
040000A6
15000000
A86B0000
A8830000
8462FFEC
D4011800
8462FFF0
D4011804
D4012008
18600001
A8631B7F
0400092F
15000000
8462FFF0
9C630001
D7E21FF0
8482FFF0
8462FFE4
E4841800
13FFFFCF
15000000
A8220000
8441FFF8
8521FFFC
85C1FFF4
44004800
15000000
D7E117F8
9C410000
D7E14FFC
9C21FFE8
D7E21FEC
9C600000
D7E21FF4
0000000F
15000000
8462FFF4
84630000
D7E21FF0
8482FFF0
8462FFEC
E4241800
10000004
15000000
0000000B
15000000
8462FFF4
9C630004
D7E21FF4
8462FFF4
188003FF
A884FFFF
E4A32000
13FFFFEF
15000000
8462FFF4
D4011800
18600001
A8631BB4
040008FF
15000000
8462FFF4
A9630000
A8220000
8441FFF8
8521FFFC
44004800
15000000
D7E117F8
9C410000
D7E14FFC
9C21FFE8
18609500
A8630200
94630000
A463FFFF
D7E21FF4
8462FFF4
04000832
15000000
E06B0004
E08C0004
18A00001
A8A51BF0
84C50004
84A50000
04000349
15000000
E06B0004
E08C0004
18A00001
A8A51BF8
84C50004
84A50000
04000050
15000000
E06B0004
E08C0004
18A00001
A8A51C00
84C50004
84A50000
04000534
15000000
E06B0004
E08C0004
D4011800
D4012004
8462FFF4
D4011808
18600001
A8631BC3
040008CA
15000000
8462FFF4
A9630000
A8220000
8441FFF8
8521FFFC
44004800
15000000
D7E117FC
9C410000
9C21FFF4
D7E21FF4
8462FFF4
B8630044
D7E21FF8
18609600
A8630004
8482FFF8
A484FFFF
DC032000
A8220000
8441FFFC
44004800
15000000
D7E117F8
9C410000
D7E14FFC
9C21FFF0
D7E21FF4
D7E227F0
18609100
A8632004
9C80AAAA
DC032000
18609100
A8632000
9C80AAAA
DC032000
18600001
A8631C08
040008E7
15000000
18600220
18800221
07FFFE76
15000000
9C600000
A9630000
A8220000
8441FFF8
8521FFFC
44004800
15000000
9C21FFFC
D4014800
04000808
15000000
9D670000
85210000
44004800
9C210004
D7E1C7EC
BB030054
D7E1F7F8
BBC3005F
D7E117D8
D7E177DC
D7E197E0
D7E1B7E8
D7E1D7F0
D7E1E7F4
D7E14FFC
D7E10FD4
D7E1A7E4
A71807FF
9C21FFC4
1840000F
BC180000
A842FFFF
D401F004
AA440000
AB450000
AB860000
AAC40000
10000045
E1C31003
BC1807FF
10000028
E24E2004
18600010
B844005D
E1CE1804
9E800000
B9CE0003
BAC40003
9F18FC01
E1CE1004
D401A000
BA5A0054
1860000F
A8BC0000
A65207FF
A863FFFF
BC120000
E05A1803
1000004E
BB5A005F
BC1207FF
10000043
18800010
B97C005D
E0422004
B8BC0003
B8420003
9E52FC01
9CC00000
E0425804
E066A004
18E00001
B8630002
A8E71C18
E09AF005
E0633800
AB840000
84630000
44001800
E2589002
BC120000
0C000054
9C400003
9C400002
A9D20000
9E800008
AAD20000
03FFFFDC
D4011000
A9C20000
AAC50000
D401D004
D4013000
84410000
BC020002
10000049
87810004
BC020003
10000295
BC020001
0C000246
9C400000
84810004
A9C20000
00000044
AAC20000
E04E2004
BC020000
10000034
9C400001
BC0E0000
100001E8
15000000
040007DE
A86E0000
A88B0000
9CA00028
9EC4FFF8
E0A52002
E1CEB008
E0B22848
E2D2B008
E1C57004
9E800000
9F00FC0D
D401A000
03FFFFB5
E3182002
E382E004
BC1C0000
0FFFFFC4
9CC00003
A85C0000
9CC00002
03FFFFC0
A8BC0000
E062E004
BC030000
10000013
A8B20000
BC020000
100001C1
15000000
040007C0
A8620000
A86B0000
9C800028
9CA3FFF8
E0841802
E0422808
E09C2048
E0BC2808
E0441004
9E40FC0D
9CC00000
03FFFFAB
E2521802
A8520000
03FFFFA8
9CC00001
9E800004
A9D80000
AAD80000
03FFFF90
D4011000
9E80000C
03FFFF8D
D4011000
9DC00000
A49C0001
9C4007FF
AACE0000
18A0000F
B8420014
A8A5FFFF
B884001F
E1CE2803
9C21003C
E1CE1004
A8760000
E1CE2004
8521FFFC
A84E0000
8421FFD4
E1620004
E1830004
85C1FFDC
8441FFD8
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
19C0000F
9C800000
A9CEFFFF
9EC0FFFF
03FFFFE4
9C4007FF
9C400000
A9C20000
03FFFFE0
AAC20000
18800008
E06E2003
BC230000
1000018F
18E00008
18A0000F
E1CE2004
A8A5FFFF
A89E0000
E1CE2803
03FFFFD4
9C4007FF
E44E1000
10000012
B8960041
E4762800
0C00019B
9C600001
A46300FF
BC030000
10000007
E06E1005
E0801802
E0641804
BD830000
0C000006
B8960041
D401B008
9E52FFFF
00000007
9EC00000
B86E001F
BAD6001F
B9CE0041
E0641804
D4011808
BB050058
B8420008
A86E0000
BA850008
E3181004
BB580050
A458FFFF
A89A0000
04000716
D4011000
A86E0000
E1CB1306
A89A0000
07FFFF07
ABCB0000
84610008
B96B0010
B8430050
E04B1004
E4AE1000
10000013
15000000
E042C000
E4B81000
0C000166
9C600001
A46300FF
BC030000
1000017F
E44E1000
10000003
9C600001
9C600000
A46300FF
BC230000
0C000178
15000000
9FDEFFFE
E042C000
E0427002
A89A0000
040006F5
A8620000
A8620000
84410000
A89A0000
E04B1306
A9CB0000
07FFFEE4
D4011004
84610008
B96B0010
A443FFFF
E16B1004
84410004
E4A25800
10000014
15000000
E16BC000
E4B85800
0C000140
9C400001
A44200FF
BC020000
10000159
84410004
E4425800
10000003
9C400001
9C400000
A44200FF
BC220000
0C000151
15000000
9DCEFFFE
E16BC000
B87E0010
A454FFFF
BBD40050
E0EE1804
84610004
A487FFFF
B8A70050
E0C41306
E1051306
E16B1802
E064F306
B8860050
E0681800
E0632000
E4A81800
10000004
E0A5F306
18800001
E0A52000
B8830050
B8630010
A4C6FFFF
E0A52000
E48B2800
1000000F
E0633000
E08B2805
E0C02002
E0862004
BD840000
10000133
E4961800
10000003
9C800001
9C800000
A48400FF
BC040000
1000002F
A9C70000
E2D6A000
9DC7FFFF
E496A000
0C000104
9C800001
E084C000
E16B2000
E4985800
1000000F
E4455800
E08BC005
E0C02002
E0862004
BD840000
1000001F
E4B4B000
10000003
9C800001
9C800000
A48400FF
BC040000
10000018
E4455800
1000000F
15000000
E0855805
E0C02002
E0862004
BD840000
10000010
E443B000
10000003
9C800001
9C800000
A48400FF
BC040000
10000009
15000000
E2D6A000
9DC7FFFE
E496A000
0C0000ED
9C800001
E084C000
E16B2000
E0761802
E16B2802
E443B000
D4011804
10000003
9EC00001
9EC00000
E2CBB002
E416C000
1000010D
A8760000
04000673
A89A0000
84A10000
A8760000
E2CB2B06
A89A0000
07FFFE63
D4015808
84E10004
B96B0010
B8670050
E16B1804
E4B65800
10000015
15000000
E16BC000
E4B85800
10000003
9C600001
9C600000
A46300FF
BC030000
1000011D
E4565800
10000003
9C600001
9C600000
A46300FF
BC230000
0C000116
84810008
E16BC000
9C84FFFE
D4012008
E2CBB002
A89A0000
0400064F
A8760000
84A10000
A8760000
E2CB2B06
A89A0000
07FFFE3F
D401580C
84E10004
B96B0010
A467FFFF
E16B1804
E4B65800
10000016
84A10008
E16BC000
E4B85800
10000003
9C600001
9C600000
A46300FF
BC030000
100000FD
E4565800
10000003
9C600001
9C600000
A46300FF
BC230000
0C0000F6
8481000C
E16BC000
9C84FFFE
D401200C
84A10008
84E1000C
B8C50010
E16BB002
E0C73004
B8E60050
A486FFFF
E0641306
E0471306
E084F306
B8A30050
E0822000
E0842800
E4A22000
10000004
E3C7F306
18400001
E3DE1000
B8A40050
B8440010
A463FFFF
E3DE2800
E48BF000
1000000D
E0421800
E08BF005
E0601002
E0A02002
E0631004
E0A52004
BD850000
1000008F
B863005F
BC030000
1000008C
15000000
E16BC000
E4B85800
10000030
9EC6FFFF
E2941005
E08BF005
E040A002
E282A004
B874005F
E0402002
E0822004
BD840000
10000093
BC030000
0C000091
15000000
9C5203FF
BDA20000
10000083
A4760007
BC030000
1000000D
18800100
A476000F
BC030004
10000009
9C760004
E483B000
10000003
9C800001
9C800000
E1CE2000
AAC30000
18800100
E06E2003
BC030000
10000007
BDA207FE
18A0FEFF
9C520400
A8A5FFFF
E1CE2803
BDA207FE
10000061
B86E001D
9EC00000
A49C0001
9C4007FF
03FFFE75
A9D60000
E45E5800
10000044
E074A000
E09E5805
E0602002
E0632004
BD830000
10000009
E4941000
10000003
9C600001
9C600000
A46300FF
BC230000
10000036
15000000
E0541005
E0601002
E0431004
03FFFFC4
B862005F
04000601
A87C0000
9C6B0020
BD430027
0FFFFE40
9D6BFFF8
A8B20000
03FFFE44
E05C5808
040005F8
A8640000
9C8B0020
BD440027
0FFFFE19
9D6BFFF8
AAD80000
03FFFE1D
E1D25808
E0623803
BC230000
10000010
18600008
E1C23804
1840000F
A89A0000
A842FFFF
AAC50000
E1CE1003
03FFFE42
9C4007FF
03FFFEFE
9C800000
03FFFEC2
9C400000
03FFFE9C
9C600000
18A0000F
E1CE1804
A8A5FFFF
A89E0000
E1CE2803
03FFFE35
9C4007FF
03FFFE67
9C600000
03FFFF15
9C800000
E074A000
9EC6FFFE
E483A000
10000003
9C800001
9C800000
E0421805
E304C000
E0601002
E16BC000
E0431004
E08BF005
03FFFF87
B862005F
03FFFEB3
9DCEFFFF
03FFFE8C
9FDEFFFF
03FFFF03
A9C70000
03FFFF7F
AAC60000
18E0000F
BAD60043
B9CE0043
A8E7FFFF
A44207FF
E2C3B004
E1CE3803
03FFFE12
A49C0001
9C40FC02
E0429002
BDA20038
1000000D
BD42001F
9C400000
A49C0001
A9C20000
03FFFE08
AAC20000
03FFFF71
AAD60001
03FFFF6F
9EC0FFFF
03FFFF6D
87810004
1000002C
BC020020
9E52041E
E0961048
E2D69008
E24E9008
E060B002
E0849004
E2C3B004
B876005F
E0841804
A4640007
BC230000
0C00000D
E04E1048
A464000F
BC030004
10000009
15000000
9C640004
E4832000
10000003
9CA00001
9CA00000
E0422800
A8830000
18A00080
E0622803
BC030000
10000023
18E0000F
9DC00000
A49C0001
9C400001
03FFFDDE
AACE0000
84610008
9C63FFFF
03FFFEED
D4011808
8461000C
9C63FFFF
03FFFF0D
D401180C
9C40FBE2
E0429002
1000001B
E04E1048
9E52043E
E1CE9008
E2CEB004
E080B002
E084B004
B884005F
E0841004
A4640007
BC230000
0C00000B
A9C30000
A464000F
BC230004
13FFFFD6
9C400000
18E0000F
B9C20043
A8E7FFFF
B862001D
E1CE3803
BAC40043
9C400000
A49C0001
03FFFDB9
E2D61804
03FFFFE9
9DC00000
18400008
1860000F
E1CE1004
A863FFFF
84810004
E1CE1803
03FFFDAF
9C4007FF
D7E1C7EC
BB030054
D7E1B7E8
BAC3005F
D7E117D8
D7E197E0
D7E1D7F0
D7E1E7F4
D7E1F7F8
D7E14FFC
D7E10FD4
D7E177DC
D7E1A7E4
AB440000
9C21FFCC
A71807FF
AA440000
1880000F
BC180000
A884FFFF
D401B004
ABC50000
AB860000
10000056
E0432003
BC1807FF
10000027
18A00010
B87A005D
E0422804
9E800000
B8420003
BA5A0003
9F18FC01
E0421804
D401A000
B9DE0054
18A0000F
A87C0000
A5CE07FF
A8A5FFFF
BC0E0000
E35E2803
10000060
BBDE005F
BC0E07FF
10000055
19600010
B87C0003
E35A5804
B97C005D
BB5A0003
9DCEFC01
9C800000
E35A5804
E284A004
18A00001
BA940002
A8A51C58
E1D87000
E2942800
E0DEB005
84B40000
44002800
9CEE0001
E342D004
BC1A0000
0C00006E
9D600003
9C800002
A85A0000
9E800008
AA5A0000
03FFFFDB
D4012000
D4013004
84A10000
BC050002
0C000052
BC050003
84410004
9E400000
A6C20001
9F4007FF
A8520000
1960000F
BB5A0014
A96BFFFF
BAD6001F
E0425803
9C210034
E042D004
A8B20000
E042B004
8521FFFC
A8820000
8421FFD4
E1640004
E1850004
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
E062D004
BC030000
1000003D
9C600001
BC020000
1000010B
15000000
040004DC
A8620000
A88B0000
9CA00028
9E44FFF8
E0A52002
E0429008
E0BA2848
E25A9008
E0451004
9E800000
9F00FC0D
D401A000
03FFFFA3
E3182002
E39AE004
BC1C0000
0FFFFFB2
9C800003
AB5C0000
9C800002
03FFFFAE
A87C0000
E07AE004
BC030000
1000001C
A86E0000
BC1A0000
100000E4
15000000
040004BE
A87A0000
A8AB0000
9C800028
9C65FFF8
E0842802
E35A1808
E09C2048
E07C1808
E344D004
9DC0FC0D
9C800000
03FFFF99
E1CE2802
10000152
BC050001
0C000109
9F400000
84410004
AA5A0000
A6C20001
03FFFFAE
A85A0000
AB4E0000
03FFFF8D
9C800001
9E800004
A8580000
AA580000
03FFFF75
D4011800
9E80000C
03FFFF72
D4015800
1840000F
9EC00000
A842FFFF
9E40FFFF
03FFFF9D
9F4007FF
A85A0000
AA430000
D401F004
03FFFF8F
D4012000
A85A0000
AA430000
D4013004
03FFFF8A
D4012000
BA720050
BA230050
A652FFFF
A463FFFF
E0B19306
E1639306
E0839B06
B90B0050
E0A42800
E0A54000
E4A42800
10000004
E1F19B06
18800001
E1EF2000
BA9A0050
A75AFFFF
B8850010
E11A9306
E19A9B06
E2549306
B9A80050
E24C9000
A56BFFFF
E2526800
B8A50050
E4AC9000
E1A45800
10000004
E0949B06
19600001
E0845800
BA620050
A442FFFF
BAB20010
E1631306
E1911306
E0639B06
BACB0050
E1836000
A508FFFF
E18CB000
BA520050
E2B54000
E4A36000
E2449000
E0B52800
10000004
E2319B06
18600001
E2311800
E09A1306
E35A9B06
E0541306
B8640050
E05A1000
B90C0050
E0421800
B98C0010
A46BFFFF
E4BA1000
E2314000
E16C1800
10000004
E2949B06
18600001
E2941800
E1057800
E4554000
10000003
9CA00001
9CA00000
B8620010
A484FFFF
E1885800
E0632000
E44B6000
E0639000
9C800001
10000003
E1032800
9C800000
E1714000
E4454000
E1EB2000
10000003
9CA00001
9CA00000
E4521800
10000003
9C600001
9C600000
E0651804
B8420050
A46300FF
E4447800
E0A31000
10000003
9D000001
9D000000
E4515800
10000003
9C600001
9C600000
E0681804
B88C0009
A50300FF
B84F0057
E0A54000
E0846804
E0A5A000
E2402002
B8A50009
E0922004
B90C0057
E0451004
18A00100
B884005F
E0622803
BA4F0009
E0844004
BC030000
10000009
E2449004
B8920041
A6520001
B862001F
E2522004
B8420041
E2521804
A9C70000
9F4E03FF
BDBA0000
10000058
A4720007
BC030000
1000000D
18800100
A472000F
BC030004
10000009
9C720004
E4839000
10000003
9C800001
9C800000
E0422000
AA430000
18800100
E0622003
BC030000
10000007
BDBA07FE
18A0FEFF
9F4E0400
A8A5FFFF
E0422803
BDBA07FE
10000024
1960000F
9E400000
A6C60001
9F4007FF
03FFFEEF
A8520000
19600008
E0825803
BC240000
10000023
18A00008
1860000F
E0425804
A863FFFF
9F4007FF
03FFFEE3
E0421803
040003DC
A87C0000
9CAB0020
BD450027
0FFFFF1D
9D6BFFF8
A86E0000
03FFFF21
E35C5808
040003D3
A87A0000
9C8B0020
BD440027
0FFFFEF6
9D6BFFF8
AA580000
03FFFEFA
E05A5808
B862001D
BA520043
B8420043
A96BFFFF
A75A07FF
E2439004
E0425803
03FFFEC8
A6C60001
E09A2803
BC240000
1000000A
1880000F
1960000F
E05A2804
A96BFFFF
AADE0000
E0425803
AA430000
03FFFEBC
9F4007FF
18600008
E0421804
A884FFFF
9F4007FF
03FFFEB6
E0422003
9C60FC02
E0637002
BDA30038
1000000A
BD43001F
9F400000
A6C60001
A85A0000
03FFFEAC
AA5A0000
A9C70000
03FFFF9B
84C10004
10000025
9C80FBE2
9DCE041E
E0921848
E2527008
E0621848
E1C27008
E0409002
E2429004
E0847004
B852005F
E0841004
A4440007
BC220000
0C00000E
18A00080
A444000F
BC020004
1000000B
E0432803
9C440004
E4822000
10000003
9CA00001
9CA00000
E0632800
A8820000
18A00080
E0432803
BC020000
1000001B
1960000F
9C400000
A6C60001
9F400001
03FFFE85
AA420000
BC030020
E0847002
1000001B
E0822048
9DCE043E
E0427008
E2429004
E0409002
E2429004
B852005F
E0822004
A4640007
BC230000
0C00000B
A8430000
A444000F
BC220004
13FFFFDE
9C600000
1960000F
B8430043
A96BFFFF
B863001D
E0425803
B8840043
A6C60001
9F400000
03FFFE67
E2441804
03FFFFE9
9C400000
18600008
18A0000F
E0421804
84810004
A8A5FFFF
A6C40001
E0422803
03FFFE5C
9F4007FF
D7E117EC
1840000F
B9850054
A842FFFF
D7E177F0
E0E31003
E1051003
A58C07FF
B9C30054
B9670003
B9A6005D
B863005F
B8E4005D
B9080003
D7E197F4
D7E14FFC
D7E10FE8
D7E1A7F8
BC2C07FF
9C21FFE8
A5CE07FF
AA430000
E0EB3804
B8440003
B8A5005F
E1086804
0C000044
B8C60003
ACA50001
E4232800
0C000046
E08E6002
E06E6002
BDA30000
100000F2
BC2C0000
1000006A
BC0E07FF
E0883004
BC040000
0C0000D1
9C63FFFF
A4620007
BC230000
0C0000BE
18600080
A462000F
BC230004
0C0000FD
9CA20004
E4851000
0C0000C4
9C600001
E0E71800
19600080
A4720001
E0875803
A8450000
BC040000
100000A4
9CAE0001
BC0507FF
100000F3
1880FF7F
1960000F
A884FFFF
B8420043
E0E72003
A96BFFFF
B887001D
B8E70043
A4A507FF
E0441004
E0E75803
1980000F
A4A507FF
A98CFFFF
B8A50014
E0E76003
B863001F
E0E72804
9C210018
E0E71804
A8A20000
A8870000
8521FFFC
8421FFE8
E1640004
E1850004
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
E0883004
BC040000
13FFFFBC
E4232800
13FFFFBE
E08E6002
BDA40000
100000E6
BC2C0000
0C00009D
BC0E07FF
13FFFFC1
BD440038
19800080
E1086004
0C00013C
BD44001F
E0C83004
9C800000
E0A03002
E0C53004
B8A6005F
E0A51000
E0E43800
E4851000
10000003
9C400001
9C400000
E0E71000
A8450000
19600080
E0875803
BC040000
1000005B
15000000
9DCE0001
BC0E07FF
100001A9
1980FF7F
B8620041
A98CFFFF
A4420001
E0E76003
E0431004
B887001F
B8E70041
03FFFF9E
E0422004
13FFFF9C
18800080
E1082004
BD430038
100000B3
BD43001F
100000DE
9C83FFE0
9CA00020
E0861848
E0A51802
E0681848
E0C62808
E1082808
E0A03002
E1082004
E0C53004
B8C6005F
E0883004
E0822002
E0E71802
E4441000
10000003
9C400001
9C400000
E0E71002
A8440000
18800080
E0672003
BC030000
1000002F
A4620007
18A0007F
A8A5FFFF
E2872803
BC140000
10000082
15000000
040002A1
A8740000
9CABFFF8
BD45001F
10000083
15000000
9C600028
E2942808
E1635802
E54E2800
E1625848
E0422808
10000080
E16BA004
E0A57002
9CE50001
BD47001F
1000009F
9C65FFE1
9DC0001F
E0623848
E0AE2802
E0EB3848
E0822808
E16B2808
9DC00000
E0402002
E1635804
E0422004
B842005F
03FFFF58
E04B1004
E0E32004
BC070000
10000209
15000000
A8E30000
A8440000
A4620007
BC230000
13FFFF53
A462000F
A4720001
B887001D
B8420043
BC0E07FF
B8E70043
1000000A
E0441004
1980000F
A4AE07FF
A98CFFFF
03FFFF62
E0E76003
E0871803
03FFFF4F
A4720001
E0823804
BC040000
100001A0
1960000F
18800008
E0E72004
A96BFFFF
A8AE0000
03FFFF55
E0E75803
03FFFF3E
9C600000
BC230000
10000066
BC0E07FF
E0C23002
E0E74002
E4461000
0C0000B8
9C400001
E0E71002
03FFFFA7
A8460000
E0A83004
BC050000
13FFFF24
9C84FFFF
BC240000
100000C2
BC0E07FF
E0C61000
E0E83800
E4861000
10000003
9C400001
A84C0000
E0E71000
03FFFF6A
A8460000
BC030000
0C00006A
9C8E0001
A48407FF
BD440001
0C0000D3
E0823002
E2874002
E4441000
10000003
9D600001
A9630000
E2945802
19800080
E0746003
BC030000
1000007D
E0E83802
E0461002
E4423000
0C0000A1
9C800001
E2872002
03FFFF86
AA450000
18A00080
A4720001
03FFFF0B
E0872803
9CE00000
03FFFF18
A8470000
04000221
A8620000
9D6B0020
9CABFFF8
BD45001F
0FFFFF81
15000000
9D6BFFD8
E54E2800
E1625808
0FFFFF84
9C400000
1980FF7F
E1CE2802
A98CFFFF
03FFFEE7
E0EB6003
E0C83004
9C600000
E0803002
E0C43004
03FFFF58
B886005F
BC040000
0C0000C2
9CAE0001
A56507FF
BD4B0001
0C000083
BC0507FF
100000E3
E0C61000
E0E83800
E4861000
10000003
9D600001
A9640000
E0E75800
B8C60041
B847001F
A9C50000
B8E70041
03FFFECC
E0423004
0FFFFF32
BD430038
03FFFEC9
A4620007
BC070020
1000006A
E06B1848
9DC0003F
E0AE2802
E16B2808
E04B1004
9CE00000
E0801002
A9C70000
E0441004
B842005F
03FFFF6A
E0421804
BC030020
1000005E
E0A82048
9C800040
E0641802
E1081808
E0C83004
9C600000
E0803002
E0C43004
B886005F
03FFFF24
E0842804
BC2E0000
0C000039
E0871004
BC0C07FF
10000086
19600080
E0601802
E0E75804
BD430038
100000A7
BD43001F
10000124
9C83FFE0
9D600020
E1A21848
E16B1802
E0671848
E0825808
E0E75808
E0402002
E0E76804
E0422004
B842005F
E0471004
E0461002
E0681802
E4423000
10000003
9CE00001
9CE00000
E0E33802
A9CC0000
03FFFF0A
AA450000
E0F42004
BC070000
0FFFFF0E
A8440000
A8670000
A8470000
03FFFF38
A9C70000
10000051
BC040020
9D600020
E0A62048
E16B2002
E0882048
E0C65808
E1085808
E1603002
E1082804
E0CB3004
B8C6005F
03FFFEBF
E0A83004
03FFFF4A
A84C0000
BC040000
1000004F
AC63FFFF
BC230000
1000004A
BC0C07FF
E0461002
E0E83802
E4423000
10000003
9C800001
A88E0000
E0E72002
A9CC0000
03FFFEE2
AA450000
03FFFF61
9C800000
0FFFFEA2
BD440038
03FFFE5E
A4620007
03FFFF9B
9D600000
03FFFFA7
9D000000
BC2E0000
100000BF
E0671004
BC030000
100000F2
E0683004
BC030000
13FFFE50
E0861000
E0E83800
E4841000
10000003
9C400001
A84E0000
E0E71000
19600080
E0475803
BC020000
100000FD
1980FF7F
A8440000
A98CFFFF
9DC00001
03FFFE40
E0E76003
BC2E0000
10000035
E0671004
BC230000
10000067
E0683004
E0483004
BC020000
100000CC
A86E0000
A8E80000
A8460000
03FFFE32
AA450000
9CA4FFE0
100000B1
E1682848
9CA00040
E0852002
E1082008
E0C83004
9C800000
E0A03002
E0C53004
B8A6005F
03FFFE6F
E0A55804
0FFFFF81
BD430038
A8E80000
A8460000
A9CC0000
03FFFE1E
AA450000
BC2E0000
1000002A
BC0C07FF
E0A71004
BC050000
10000078
15000000
AC84FFFF
BC240000
10000072
BC0C07FF
E0423000
E0E83800
E4823000
10000003
9C800001
A88E0000
E0E72000
03FFFE5C
A9CC0000
BC230000
1000004B
E0683004
BC030000
10000095
AA450000
A8E80000
A8460000
03FFFE00
9DC007FF
9CE00000
03FFFEB2
A8470000
E0471004
9C600000
E0801002
E0441004
03FFFF64
B842005F
A8E40000
A9C50000
03FFFEA8
A8440000
10000052
15000000
18A00080
E0802002
E0E72804
BD440038
10000084
BD44001F
1000008F
9CA4FFE0
9D600020
E1A22048
E16B2002
E0872048
E0A25808
E0E75808
E0402802
E0E76804
E0422804
B842005F
E0471004
E0423000
E1044000
E4823000
10000003
9CE00001
9CE00000
E0E83800
03FFFE27
A9CC0000
BC030000
13FFFDD3
A4620007
E0823002
E0674002
E4441000
10000003
9D600001
A96E0000
E0635802
19800080
E1636003
BC0B0000
13FFFE70
E0461002
E0E83802
E4423000
10000003
9C800001
9C800000
E0E72002
03FFFDBE
AA450000
BC030000
13FFFDBB
9DC007FF
B8870043
19600008
B8420043
E0645803
B8E7001D
BC030000
1000000C
E0471004
B8E80043
E0675803
BC230000
10000007
15000000
B8C60043
B848001D
A8870000
AA450000
E0423004
B8E2005D
B8840003
B8420003
9DC007FF
03FFFDA3
E0E72004
0FFFFFB6
BD440038
A8E80000
A8460000
03FFFD9D
A9CC0000
A8E40000
A8AE0000
03FFFDB9
A8440000
BC030000
10000038
E0683004
BC030000
13FFFD93
9DC007FF
B8870043
18A00008
B8420043
E0642803
B8E7001D
BC030000
13FFFFE4
E0471004
B8A80043
18E00008
E0653803
BC230000
13FFFFDE
15000000
B8C60043
B848001D
A8850000
03FFFFD9
E0423004
03FFFF54
9D000000
BC030020
1000002E
E0872048
9D600040
E06B1802
E0E71808
E0471004
9C600000
E0E01002
E0471004
B842005F
03FFFEDE
E0422004
18E0007F
9C40FFF8
A8E7FFFF
03FFFE21
9DC007FF
A8EE0000
03FFFE1E
A84E0000
E0471004
9C800000
E0A01002
E0451004
03FFFF87
B842005F
A8E80000
03FFFD60
A8460000
A8E80000
A8460000
03FFFD5C
9DC007FF
BC040020
10000013
E0A72848
9D600040
E08B2002
E0E72008
E0471004
9C800000
E0E01002
E0471004
B842005F
03FFFF73
E0422804
03FFFFD7
9CE00000
A8670000
03FFFDFF
A8470000
03FFFDF8
A8440000
03FFFFF2
9CE00000
D7E117F8
D7E14FFC
D7E10FF4
BC030000
9C21FFF4
10000012
A8430000
04000068
15000000
9C80041E
BD4B000A
1000001D
E0845802
9C60000B
9CAB0015
E1635802
1860000F
E1625848
A863FFFF
A48407FF
E0422808
00000004
E16B1803
A8830000
A9630000
1860000F
A48407FF
A863FFFF
B8840014
E16B1803
9C21000C
E08B2004
A8E20000
A8C40000
8521FFFC
8421FFF4
E1660004
E1870004
44004800
8441FFF8
9D6BFFF5
1860000F
E1625808
A863FFFF
A48407FF
9C400000
03FFFFEB
E16B1803
9C21FFFC
D4014800
9D600000
9D040000
9CA30000
E4285800
0C000036
9CE00000
E4482800
10000032
E4082800
1000002E
E48B4000
0C00000D
9DA00020
19208000
9CC0FFFF
E0654803
B8870001
9DE50000
B863005F
E1AD3000
E0E41804
E4874000
13FFFFF9
B8A50001
B8E70041
9DAD0001
9D200000
E4896800
0C00001E
9CAF0000
19E08000
9E200000
E0657803
B8870001
B863005F
E0E41804
E0C74002
E0667803
B863005F
9C800000
E4232000
10000003
B86B0001
9C800001
B8A50001
E4248800
0C000003
E1632004
9CE60000
9D290001
E4896800
13FFFFED
15000000
00000005
15000000
00000003
9D600001
9CE50000
85210000
44004800
9C210004
D7E117FC
A840FFFF
D7E10FF8
E4431000
10000011
9C21FFF8
BCA300FF
10000019
9C800000
9C800008
9D600018
18400001
E0632048
A8421C98
9C210008
E0631000
8421FFF8
8C630000
8441FFFC
44004800
E16B1802
184000FF
A842FFFF
E4A31000
0C000005
15000000
9C800010
03FFFFF0
A9640000
9C800018
03FFFFED
9D600008
03FFFFEB
9D600020
A8830000
9C600000
D7E14FFC
D7E10FF8
A8A30000
9C21FFF8
040009A9
A8C30000
9C210008
8521FFFC
44004800
8421FFF8
D7E117F8
D7E14FFC
D7E10FF4
9C800000
9C21FFF4
040009EE
A8430000
18600001
A8631D98
84630000
8483003C
BC040000
10000004
15000000
48002000
15000000
04002AA3
A8620000
D7E14FFC
D7E10FF8
9C21FFF8
A8A40000
9CC10008
0400009C
84830008
9C210008
8521FFFC
44004800
8421FFF8
D7E14FFC
D7E117F8
D7E10FF4
9C21FFF4
04001718
A8430000
A8A20000
9CC1000C
A86B0000
0400008D
848B0008
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E117F4
D7E177F8
A8440000
A9C30000
D7E14FFC
A8640000
D7E10FF0
0400003D
9C21FFD4
D401100C
18400001
9C8B0001
A8421D9E
846E0038
D4011014
9C400001
D4015810
D4011018
9C41000C
D4012008
D4011000
9C400002
BC230000
D4011004
0C00001A
844E0008
9862000C
A4832000
BC240000
10000007
9CA0DFFF
84820064
A8632000
E0842803
DC02180C
D4022064
A86E0000
A8820000
0400150A
A8A10000
BC2B0000
10000003
9D60FFFF
9D60000A
9C21002C
8521FFFC
8421FFF0
8441FFF4
44004800
85C1FFF8
040013A3
A86E0000
03FFFFE7
9862000C
D7E14FFC
D7E117F8
D7E10FF4
9C21FFF4
040016D2
A8430000
A8820000
07FFFFC3
A86B0000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
A4830003
D7E10FF8
D7E117FC
BC040000
1000003A
9C21FFF8
90A30000
BC050000
10000038
A8830000
00000007
9C840001
90A40000
BC250000
0C00002C
E1641802
9C840001
A4A40003
BC250000
13FFFFF9
15000000
1840FEFE
84A40000
A842FEFF
E0C51000
ACA5FFFF
18408080
E0A62803
A8428080
E0A51003
BC250000
10000010
15000000
9C840004
1840FEFE
84A40000
A842FEFF
E0C51000
ACA5FFFF
18408080
E0A62803
A8428080
E0A51003
BC050000
13FFFFF6
9C840004
9C84FFFC
90A40000
BC050000
10000009
E1641802
9C840001
90A40000
BC250000
13FFFFFE
9C840001
9C84FFFF
E1641802
9C210008
8421FFF8
44004800
8441FFFC
03FFFFD7
A8830000
03FFFFFA
A9650000
D7E14FFC
D7E1A7E4
D7E1D7F0
D7E10FD4
D7E117D8
D7E177DC
D7E197E0
D7E1B7E8
D7E1C7EC
D7E1E7F4
D7E1F7F8
9C21FEE4
AA830000
AB440000
D4012818
040016B9
D4013024
856B0000
A86B0000
07FFFFAB
D4015844
BC140000
10000006
D4015850
84540038
BC220000
0C0000BC
15000000
987A000C
A443FFFF
A4822000
BC240000
10000008
9CA0DFFF
849A0064
A8432000
E0642803
DC1A100C
D41A1864
A442FFFF
A4620008
BC030000
10000072
A8740000
847A0010
BC230000
0C00006D
A442001A
BC22000A
0C000075
9C400000
9EC100B0
D401102C
9C4100AF
9C600000
D4011008
9C41007C
D401B07C
D4011010
9C41006C
D4011884
D401100C
84410008
D4011880
E0561002
D4011848
D401184C
AB960000
D4011858
D4011854
D4011830
D401105C
84610018
90430000
AC620025
A46300FF
BC030000
1000008D
15000000
A44200FF
BC020000
10000089
15000000
00000005
84410018
BC230000
0C00000A
84810018
9C420001
90620000
AC830025
A48400FF
BC040000
0FFFFFF8
A46300FF
84810018
E1C22002
BC0E0000
10000010
84810084
84610080
E0847000
9C630001
84A10018
D41C7004
D41C2800
D4012084
BD430007
10000053
D4011880
9F9C0008
84E10030
E0E77000
D4013830
90620000
BC030000
10000054
9CA00000
9C600000
9C80FFFF
9C420001
D8011861
D4012014
D4012828
ABC50000
90C20000
9C820001
9C46FFE0
BC420058
10000213
18E00001
B8420002
A8E71DE4
E0423800
84420000
44001000
15000000
ABDE0010
03FFFFF3
A8440000
84410024
84E10024
84420000
9CE70004
D4011028
D4013824
84610028
BD630000
13FFFFE9
A8440000
E0601802
D4011828
ABDE0004
03FFFFE4
A8440000
A8740000
040007E6
A89A0000
BC0B0000
0C000012
15000000
945A000C
A442001A
BC22000A
13FFFF8F
9C400000
985A000E
BD820000
13FFFF8B
9C400000
A8740000
A89A0000
84A10018
0400079C
84C10024
00000004
9C21011C
9D60FFFF
9C21011C
8521FFFC
8421FFD4
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
A8740000
A89A0000
0400221F
9CA1007C
BC2B0000
1000000B
AB960000
03FFFFAA
84E10030
84410084
BC220000
0C000005
A8740000
A89A0000
04002213
9CA1007C
945A000C
A4420040
BC220000
13FFFFDF
85610030
03FFFFDF
9C21011C
04001279
A8740000
03FFFF45
987A000C
03FFFF98
84410018
A8440000
03FFFFA0
9CA0002B
84410024
9C600000
84420000
D4012018
D4011038
BC220000
84810024
D401303C
D8011861
0C00063C
9C440004
84610014
9C800000
BD830000
100005FE
84610038
040018D5
84A10014
BC2B0000
0C0006D4
84A10038
9CE00000
E16B2802
92410061
AC6BFFFF
D4015820
B863009F
D4013814
D4011024
E06B1803
D4013840
D401181C
BC120000
10000006
A45E0002
8441001C
9C420001
D401101C
A45E0002
BC020000
10000005
D4011034
8441001C
9C420002
D401101C
A71E0084
BC180000
0C00019F
84410084
84610028
8441001C
E1C31002
BD4E0000
0C000198
84610080
1A400001
BD4E0010
84810084
AA521F58
9C400010
10000008
A8A30000
0000001C
9C630001
9DCEFFF0
BD4E0010
0C000016
9F9C0008
9CA50001
9C840010
D41C9000
D41C1004
D4012084
BD450007
0FFFFFF6
D4012880
A8740000
A89A0000
040021B3
9CA1007C
BC2B0000
13FFFF9F
9DCEFFF0
84810084
BD4E0010
84A10080
13FFFFEE
AB960000
A8650000
9C630001
E04E2000
D41C9000
D41C7004
D4011084
BD430007
10000397
D4011880
9F9C0008
0000016C
92410061
A47E0010
D401303C
D4012018
BC030000
100000E0
84410024
84E10024
9C800001
9CE70004
D4013824
84420000
9C600000
9E400000
D8011861
84A10014
BD850000
10000004
9CE0FF7F
E3DE3803
84A10014
E0602802
E0632804
BD830000
1000029E
E0601002
E0631004
B863005F
BC030000
0C000299
BC240000
1000030A
A45E0001
BC020000
1000036E
9C600030
8441005C
D80118AF
9C6100AF
D4011020
D4011838
84410020
84610014
E5621800
10000003
15000000
A8430000
D401101C
9C400000
03FFFF8C
D4011040
BC250000
13FFFF07
A8440000
03FFFF05
9CA00020
ABDE0001
03FFFF02
A8440000
90C40000
BC06002A
10000684
9C440001
9CE6FFD0
A8820000
BCA70009
0C00000E
9C600000
E0631800
90C40000
B8430002
E0631000
E0671800
9CE6FFD0
BCA70009
13FFFFF9
9C840001
BD630000
0C00050F
15000000
03FFFEED
D4011814
ABDE0080
03FFFEE8
A8440000
D4012018
A49E0010
D401303C
BC040000
1000007C
84410024
84A10024
9C800000
9CA50004
D4012824
03FFFFAD
84420000
84A10024
D4012018
84450000
18800001
9CA50004
A8841DC1
9CE00030
9C600078
D4012824
9CA00078
D4012058
ABDE0002
D8013862
D8011863
9C800002
03FFFF9C
D401283C
9C400000
A8640000
D4011028
9CE6FFD0
E0421000
90C30000
B8620002
9C840001
E0421800
E0423800
9CE6FFD0
BCA70009
13FFFFF8
A8640000
03FFFEBD
D4011028
ABDE0010
D401303C
A47E0010
D4012018
D8012861
BC030000
1000009B
84410024
84610024
9C630004
D4011824
84420000
BD820000
100003C7
9CE0002D
92410061
03FFFF7D
9C800001
84410024
D401303C
84420000
D4012018
D4011048
84410024
84C10048
84420004
D8012861
A8820000
D401104C
A8640000
A8460000
84810024
9DC40008
E0830004
E0620004
04001FD3
15000000
84A10048
BC2B0001
8481004C
100003B1
A8450000
18E00001
A8640000
A8E71DDC
E0830004
E0620004
84A70000
84C70004
04002FE3
15000000
BD8B0000
10000574
9C40002D
92410061
18800001
8461003C
A8841DA4
BD430047
0C00049C
D4012038
9C400003
9C60FF7F
D401101C
9C400000
E3DE1803
D4011014
8441001C
D4017024
D4011020
84410014
03FFFEF4
D4011040
ABDE0008
03FFFE6F
A8440000
ABDE0010
D4012018
A49E0010
D401303C
BC040000
0FFFFF88
84410024
A47E0040
BC030000
10000410
84E10024
84420000
9CE70004
A442FFFF
03FFFF30
D4013824
ABDE0010
D401303C
A47E0010
D4012018
BC030000
0FFFFF24
84410024
A47E0040
BC030000
100003FA
84610024
84420000
9C630004
A442FFFF
D4011824
03FFFF1F
9C800001
18600001
D401303C
A8631DB0
D4012018
D4011858
A47E0010
D8012861
BC030000
10000042
84410024
84E10024
9CE70004
D4013824
84420000
A47E0001
BC030000
13FFFF0D
9C800002
BC020000
13FFFF0B
9C600000
9CA00030
84E1003C
D8012862
D8013863
03FFFF05
E3DE2004
84610024
9E400000
84430000
D4012018
9CA00000
9C800001
9C630004
9CE10088
D401303C
D401201C
D8011088
D8012861
D4011824
D4012020
D4019014
D4019040
03FFFEA9
D4013838
A47E0010
D401303C
D4012018
D8012861
BC030000
0FFFFF69
84410024
A47E0040
BC030000
100003D2
84A10024
84810024
98420002
9C840004
03FFFF64
D4012024
ABDE0040
03FFFE0E
A8440000
D8012861
18A00001
A47E0010
A8A51DC1
D401303C
D4012018
D4012858
BC030000
0FFFFFC2
84410024
A47E0040
BC030000
100003A1
84610024
84420000
9C630004
A442FFFF
03FFFFBD
D4011824
A45E0010
D4012018
BC020000
0C00001E
D8012861
A45E0040
BC020000
1000001B
84610024
84A10024
84E10030
84450000
9CA50004
DC023800
03FFFDB6
D4012824
D401303C
D4012018
BC060000
13FFFE31
D8012861
9E400000
9C400001
9C600000
9C810088
D401101C
D8013088
D8011861
D4011020
D4019014
D4019040
03FFFE62
D4012038
84610024
84810030
84430000
9C630004
D4011824
03FFFD9E
D4022000
84410084
BC120000
1000000F
84A10034
84610080
9C810061
9C630001
9C420001
D41C2000
9C800001
D4011084
D41C2004
BD430007
100001BE
D4011880
9F9C0008
84A10034
BC050000
1000000F
BC380080
84610080
9C420002
9C630001
9CE10062
9C800002
D41C3800
D41C2004
D4011084
BD430007
100001B7
D4011880
9F9C0008
BC380080
0C000153
84610028
84A10014
84E10020
E2453802
BDB20000
1000002C
84610080
19C00001
BD520010
A9CE1F48
9F000010
10000008
A8A30000
0000001C
9C630001
9E52FFF0
BD520010
0C000016
9F9C0008
9CA50001
9C420010
D41C7000
D41CC004
D4011084
BD450007
0FFFFFF6
D4012880
A8740000
A89A0000
04001FF5
9CA1007C
BC2B0000
13FFFDE1
9E52FFF0
84410084
BD520010
84A10080
13FFFFEE
AB960000
A8650000
9C630001
E0429000
D41C7000
D41C9004
D4011084
BD430007
10000172
D4011880
9F9C0008
A47E0100
BC230000
1000009F
84E1003C
84610020
84810038
E0421800
84610080
84A10020
9C630001
D41C2000
D41C2804
D4011084
BD430007
1000008A
D4011880
9F9C0008
A47E0004
BC030000
10000039
8461001C
84610028
8481001C
E1C32002
BDAE0000
10000032
84610080
1A400001
BD4E0010
AA521F58
9F000010
10000008
A8A30000
0000001C
9C630001
9DCEFFF0
BD4E0010
0C000016
9F9C0008
9CA50001
9C420010
D41C9000
D41CC004
D4011084
BD450007
0FFFFFF6
D4012880
A8740000
A89A0000
04001FB0
9CA1007C
BC2B0000
13FFFD9C
9DCEFFF0
84410084
BD4E0010
84A10080
13FFFFEE
AB960000
A8650000
9C630001
E0427000
D41C9000
D41C7004
D4011084
BDA30007
10000009
D4011880
A8740000
A89A0000
04001F9B
9CA1007C
BC2B0000
13FFFD87
84410084
8461001C
84A10028
E5632800
10000003
BC220000
A8650000
84410030
E0421800
10000110
D4011030
9C600000
AB960000
03FFFCF2
D4011880
86410080
BD470001
9E520001
0C000209
9C420001
84610038
D4011084
D41C1800
9C600001
D4019080
BD520007
10000208
D41C1804
9F9C0008
84810050
9E520001
E0422000
84A10044
D41C2004
D41C2800
D4011084
BD520007
10000207
D4019080
9F9C0008
84810048
8461004C
18E00001
A9840000
A8E71DDC
A9A30000
84A70000
84C70004
E06C0004
E08D0004
04002DA0
15000000
BC2B0000
0C000161
84E1002C
8481002C
84A10038
9C64FFFF
9C850001
9E520001
E0421800
D41C2000
D41C1804
D4011084
BD520007
100000CE
D4019080
9F9C0008
84A10054
9E520001
E0422800
9CE1006C
D41C2804
D41C3800
D4011084
BD520007
0FFFFF7A
D4019080
A8740000
A89A0000
04001F47
9CA1007C
BC2B0000
13FFFD33
84410084
03FFFF72
AB960000
BDA70065
13FFFFB7
84E1002C
84810048
8461004C
A9840000
18800001
A9A30000
A8841DDC
84A40000
84C40004
E06C0004
E08D0004
04002D6E
15000000
BC0B0000
0C0000D9
86410064
18800001
84610080
A8841DD9
9C630001
9C420001
D41C2000
9C800001
D4011084
D41C2004
BD430007
10000281
D4011880
9F9C0008
84610064
84A1002C
E5832800
10000007
84E10050
A47E0001
BC030000
13FFFF4B
A47E0004
84E10050
84610080
E0423800
9C630001
84810044
D41C3804
D41C2000
D4011084
BD430007
100002FC
D4011880
9F9C0008
84A1002C
9E45FFFF
BDB20000
13FFFF39
84610080
19C00001
BD520010
A9CE1F48
9F000010
10000009
A8A30000
00000122
9C630001
9F9C0008
9E52FFF0
BD520010
0C00011C
A8650000
9CA50001
9C420010
D41C7000
D41CC004
D4011084
BD450007
0FFFFFF5
D4012880
A8740000
A89A0000
04001EF0
9CA1007C
BC2B0000
13FFFCDC
84410084
84A10080
03FFFFEC
AB960000
BC040001
100000CF
BC040002
D401B038
0C00000F
A8960000
84A10058
A462000F
B8420044
E0651800
9C84FFFF
8C630000
BC220000
13FFFFFA
D8041800
D4012038
E0562002
03FFFD62
D4011020
A4620007
B8420043
9C84FFFF
9C630030
BC220000
13FFFFFB
D8041800
A45E0001
BC220000
0FFFFFF4
D4012038
BC230030
0C0002E9
84610038
9CA00030
9C63FFFF
DBE42FFF
E0561802
D4011838
03FFFD4D
D4011020
8481001C
E2432002
BDB20000
13FFFEAC
19C00001
84610080
BD520010
A9CE1F48
9F000010
10000008
A8A30000
0000001C
9C630001
9E52FFF0
BD520010
0C000016
9F9C0008
9CA50001
9C420010
D41C7000
D41CC004
D4011084
BD450007
0FFFFFF6
D4012880
A8740000
A89A0000
04001EA5
9CA1007C
BC2B0000
13FFFC91
9E52FFF0
84410084
BD520010
84A10080
13FFFFEE
AB960000
A8650000
9C630001
E0429000
D41C7000
D41C9004
D4011084
BD430007
10000143
D4011880
03FFFE81
9F9C0008
9E520001
E042C000
D41C7000
D41CC004
D4011084
BD520007
0FFFFF36
D4019080
A8740000
A89A0000
04001E86
9CA1007C
BC2B0000
13FFFC72
84410084
86410080
03FFFF2D
AB960000
A8740000
A89A0000
04001E7C
9CA1007C
BC2B0000
0FFFFEEE
9C600000
03FFFC67
945A000C
D4011820
03FFFCFF
D401B038
A8740000
A89A0000
04001E70
9CA1007C
BC2B0000
13FFFC5C
84410084
03FFFE8A
AB960000
A8740000
A89A0000
04001E67
9CA1007C
BC2B0000
13FFFC53
84410084
03FFFE3E
AB960000
A8740000
A89A0000
04001E5E
9CA1007C
BC2B0000
13FFFC4A
84410084
03FFFE45
AB960000
BD520000
0C0001BC
84A1002C
84610038
84E10040
E0632800
E5A53800
D4011814
10000003
A9C50000
A9C70000
BDAE0000
1000000C
84610080
E0427000
9C630001
84810038
D41C7004
D41C2000
D4011084
BD430007
10000259
D4011880
9F9C0008
AE4EFFFF
84A10040
BA52009F
E1CE9003
E2457002
BDB20000
1000006B
84610080
19C00001
BD520010
A9CE1F48
9F000010
10000009
A8A30000
00000181
9C630001
9F9C0008
9E52FFF0
BD520010
0C00017B
A8650000
9CA50001
9C420010
D41C7000
D41CC004
D4011084
BD450007
0FFFFFF5
D4012880
A8740000
A89A0000
04001E20
9CA1007C
BC2B0000
13FFFC0C
84410084
84A10080
03FFFFEC
AB960000
BC420009
100000B6
A9D60000
9C420030
8461005C
9C8100AF
D4011820
D80110AF
03FFFC9B
D4012038
D4012020
03FFFC98
D401B038
A8740000
A89A0000
04001E09
9CA1007C
BC2B0000
13FFFBF5
92410061
84410084
03FFFDD0
AB960000
9F07FFFF
BDB80000
13FFFEAC
19C00001
BDB80010
0C000009
A9CE1F48
03FFFF6B
9E520001
9F9C0008
9F18FFF0
BD580010
0FFFFF65
15000000
9E520001
9C420010
9C600010
D41C7000
D41C1804
D4011084
BD520007
0FFFFFF4
D4019080
A8740000
A89A0000
04001DE8
9CA1007C
BC2B0000
13FFFBD4
84410084
86410080
03FFFFEB
AB960000
9C630001
E0429000
D41C7000
D41C9004
D4011084
BD430007
0FFFFE09
D4011880
03FFFE90
A8740000
A8740000
A89A0000
04001DD4
9CA1007C
BC2B0000
13FFFBC0
84410084
AB960000
86410064
8481002C
84E10038
84610040
E5922000
10000040
E3071800
A47E0001
BC030000
0C00003C
15000000
8461002C
84810014
E2439002
E064C002
E5B21800
10000003
A9D20000
A9C30000
BDAE0000
1000000B
84610080
E0427000
9C630001
D41CC000
D41C7004
D4011084
BD430007
100001EA
D4011880
9F9C0008
AC6EFFFF
B863009F
E1CE1803
E2527002
BDB20000
13FFFDDA
84610080
19C00001
BD520010
A9CE1F48
9F000010
10000009
A8A30000
03FFFFC3
9C630001
9F9C0008
9E52FFF0
BD520010
0FFFFFBD
A8650000
9CA50001
9C420010
D41C7000
D41CC004
D4011084
BD450007
0FFFFFF5
D4012880
A8740000
A89A0000
04001D91
9CA1007C
BC2B0000
13FFFB7D
84410084
84A10080
03FFFFEC
AB960000
84A10050
84610080
E0422800
9C630001
84E10044
D41C2804
D41C3800
D4011084
BD430007
100001AE
D4011880
03FFFFBB
9F9C0008
A47E0001
BC030000
0FFFFDF7
84810038
9C600001
03FFFE1E
D41C2000
A8740000
A89A0000
04001D73
9CA1007C
BC2B0000
13FFFB5F
84410084
86410080
03FFFDF3
AB960000
A8740000
A89A0000
04001D69
9CA1007C
BC2B0000
13FFFB55
84410084
86410080
03FFFDF4
AB960000
A8620000
9C80000A
07FFF155
9DCEFFFF
9D6B0030
A8620000
9C80000A
07FFF95A
D80E5800
BC2B0000
13FFFFF6
A84B0000
E0567002
D4017038
03FFFBDE
D4011020
A8740000
A89A0000
04001D4F
9CA1007C
BC2B0000
13FFFB3B
84410084
03FFFD39
AB960000
E0401002
D8013861
9E40002D
03FFFBB6
9C800001
A8640000
E0830004
E0620004
04001C1A
15000000
BC2B0000
0C0000E8
18800001
84410014
8461003C
9C80FFDF
BC22FFFF
0C000103
E2432003
AC520047
E0601002
E0431004
BD820000
100000FF
84A10014
E0402802
E0422804
BD620000
0C0000FA
84410048
9E400047
BD820000
9C400001
D4011014
A85E0100
1000021E
D4011024
9C400000
87010048
D4011034
8441004C
9C610068
A8A20000
9C410074
D4011800
A8980000
D4011004
A8740000
9CC00002
84E10014
0400048B
9D010064
BC320047
10000260
D4015838
A47E0001
84E10038
84810014
BC230000
0C000219
E0472000
8461004C
18800001
A9980000
A8841DDC
A9A30000
84A40000
84C40004
E06C0004
E08D0004
04002B3D
15000000
BC0B0000
1000000E
A8620000
84610074
E4A21800
1000000B
84E10038
9C830001
9CA00030
D4012074
D8032800
84610074
E4421800
13FFFFFC
9C830001
84E10038
BC320047
E0633802
1000017D
D401182C
84410064
84810014
E5841000
10000003
9C600001
9C600000
A46300FF
BC230000
10000188
BD82FFFD
10000003
9C800001
A8830000
A48400FF
BC040000
0C000181
9C800067
D4011040
D401203C
8441002C
84610040
E5421800
100001D5
84410040
A45E0001
BC220000
100001E5
84410040
AC43FFFF
D4011820
B842009F
E0431003
84E10034
BC270000
10000121
9C60002D
87C10024
92410061
D401101C
D4017024
03FFFAE3
D4013814
84810024
9C840004
D4012024
03FFFC1E
84420000
84810024
9C840004
D4012024
9C800001
03FFFB27
84420000
84810024
9C840004
D4012024
A8830000
03FFFB21
84420000
9C630001
E0429000
D41C7000
D41C9004
D4011084
BD430007
13FFFED5
D4011880
03FFFEDB
9F9C0008
9CA50004
D4012824
03FFFB95
84420000
A8740000
A89A0000
04001CA1
9CA1007C
BC2B0000
13FFFA8D
84410084
03FFFD7B
AB960000
18800001
84610080
A8841DD9
9C630001
9C420001
D41C2000
9C800001
D4011084
D41C2004
BD430007
10000052
D4011880
9F9C0008
84E1002C
E0723804
BC230000
10000007
84610050
A47E0001
BC030000
13FFFCB7
A47E0004
84610050
84810044
E0421800
84610080
84A10050
9C630001
D41C2000
D41C2804
D4011084
BD430007
10000168
D4011880
9F9C0008
E2409002
BDB20000
10000074
19C00001
BDB20010
A9CE1F48
9F000010
0C000009
A8A30000
00000093
9C630001
9F9C0008
9E52FFF0
BD520010
0C00008D
A8650000
9CA50001
9C420010
D41C7000
D41CC004
D4011084
BD450007
0FFFFFF5
D4012880
A8740000
A89A0000
04001C5D
9CA1007C
BC2B0000
13FFFA49
84410084
84A10080
03FFFFEC
AB960000
8461003C
A8841DAC
BD430047
10000005
D4012038
18A00001
A8A51DA8
D4012838
9C400003
9C60FF7F
D401101C
9C400000
E3DE1803
D4011014
03FFFB6E
92410061
18A00001
A8A51DA0
03FFFB64
D4012838
9C60FFFF
03FFF9DF
D4011814
A8740000
A89A0000
04001C3C
9CA1007C
BC2B0000
13FFFA28
86410064
84410084
03FFFFA9
AB960000
9C400006
D4011014
84410048
BD620000
A85E0100
0C000128
D4011024
9C400000
87010048
D4011034
BC120046
10000088
8441004C
BC320045
13FFFF07
84610014
9CC10068
9C430001
8461004C
D4013000
A8A30000
9C610074
A8980000
D4011804
9CC00002
A8740000
A8E20000
0400038E
9D010064
D4015838
84810038
03FFFF0A
E0441000
A8740000
A89A0000
04001C11
9CA1007C
BC2B0000
13FFF9FD
84410084
03FFFD00
AB960000
A8740000
A89A0000
04001C08
9CA1007C
BC2B0000
13FFF9F4
84410084
84610080
AB960000
84E1002C
9C630001
E0423800
84810038
D41C3804
D41C2000
D4011084
BD430007
0FFFFC28
D4011880
03FFFCAF
A8740000
07FFF8D3
D4012014
AC6BFFFF
D4011024
B843009F
84A10014
D4015820
E04B1003
92410061
D4012840
03FFFA0A
D401101C
A8740000
A89A0000
04001BE7
9CA1007C
BC2B0000
13FFF9D3
84410084
03FFFDA3
AB960000
84410038
E0561002
03FFFA69
D4011020
9C630001
E0429000
D41C7000
D41C9004
D4011084
BD430007
13FFFFCC
D4011880
03FFFFD3
9F9C0008
A8740000
A89A0000
04001BD0
9CA1007C
BC2B0000
13FFF9BC
86410064
84410084
03FFFE07
AB960000
A8740000
A89A0000
04001BC6
9CA1007C
BC2B0000
13FFF9B2
86410064
84A1002C
84410084
E2459002
03FFFE0F
AB960000
86410014
BCB20006
10000003
15000000
9E400006
D4019020
D4011024
84A10020
18E00001
AC65FFFF
9E400000
B843009F
A8E71DD2
D4019014
E0451003
D4019040
D401101C
03FFF9D0
D4013838
D401101C
9C400000
87C10024
D8011861
D4017024
9E40002D
03FFF9C5
D4011014
9C610068
A8A20000
9C410074
D4011800
D4011004
A8980000
A8740000
9CC00003
84E10014
0400030D
9D010064
8C4B0000
84A10014
AC420030
E0AB2800
9C42FFFF
D4015838
BD620000
10000099
D401281C
8441004C
18800001
A9A20000
A9980000
A8841DDC
84A40000
84C40004
E06C0004
E08D0004
040029BF
9C400001
BC2B0000
10000004
A44200FF
A84B0000
A44200FF
BC220000
0C000086
84A10014
9C400001
E0422802
D4011064
84E1001C
03FFFE6B
E0471000
9E40002D
03FFFA8E
D8011061
84E1003C
BD470065
0C0000BE
8481003C
84410064
BC040066
0FFFFE92
D4011040
BDA20000
100000A0
84410014
BC220000
10000081
9E420001
A45E0001
BC220000
1000007B
15000000
84410040
03FFFE92
D4011020
84A1003C
9CA5FFFE
D401283C
9C42FFFF
8461003C
D4011064
BD620000
0C000097
D801186C
9CA0002B
D801286D
BDA20009
1000005E
9C800030
9F01007B
AA580000
A8620000
9C80000A
0400268D
9E52FFFF
9D6B0030
A8620000
9C80000A
0400266F
D8125800
BD4B0009
13FFFFF6
A84B0000
9C4B0030
9C72FFFF
B8420018
E463C000
B8420098
1000008C
DBF217FF
00000003
9C81006E
90430000
9C630001
D8041000
E423C000
13FFFFFC
9C840001
84E10010
9C61006E
E0479002
E0431000
84A1000C
E0422802
D4011054
8441002C
84610054
BD420001
E0421800
0C000054
D4011020
84410020
9C420001
D4011020
9C400000
84610020
D4011040
AC43FFFF
B842009F
03FFFE50
E0431003
84810014
92410061
D401201C
D4012020
D4015814
D4011024
03FFF933
D4015840
A8740000
A89A0000
04001B10
9CA1007C
BC2B0000
13FFF8FC
86410064
84410084
84610080
03FFFE92
AB960000
84410048
18608000
E3021800
9C40002D
03FFFED9
D4011034
BD420000
0C000046
9C400001
8481002C
E0422000
D4011020
AC42FFFF
84A10020
B842009F
03FFFE2C
E0451003
03FFFF7F
84410064
03FFFE03
84610074
9C420030
D801106F
D801206E
03FFFFC2
9C410070
9C420001
D4011020
AC42FFFF
84610020
B842009F
03FFFE1C
E0431003
84410014
9E420001
84410040
E2429000
AC52FFFF
D4019020
B842009F
03FFFE13
E0521003
84610024
84810024
84630000
9C840004
D4011814
BD630000
13FFF874
D4012024
9CE0FFFF
03FFF871
D4013814
A47E0001
BC230000
13FFFFAC
15000000
AC42FFFF
84810020
B842009F
D4011840
03FFFDFE
E0441003
BC220000
10000012
84410014
A45E0001
BC020000
0C00000D
15000000
9C400001
03FFFDF4
D4011020
9C80002D
E0401002
03FFFF6B
D801206D
9C400002
84610040
03FFFFBA
E0421802
84410014
03FFFFC9
9C420002
03FFFE9D
84410014
03FFFF58
84410064
03FFFF82
9C41006E
D7E14FFC
D7E117F0
D7E177F4
D7E197F8
D7E10FEC
9C21FFEC
AA430000
A9C40000
04000E4B
A8450000
A8920000
A8AE0000
A8C20000
07FFF7C0
A86B0000
9C210014
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
94E4000C
D7E117F0
D7E177F4
A8440000
85C40064
9C80FFFD
D7E197F8
E0E72003
D7E14FFC
D7E10FEC
9C21FB84
9D000400
DC01380C
94E2000E
9D610068
85A2001C
85820024
DC01380E
A8810000
9CE00000
D4017064
AA430000
D401681C
D4016024
D4015800
D4015810
D4014008
D4014014
07FFF79B
D4013818
BD8B0000
10000008
A9CB0000
A8720000
040009AD
A8810000
BC0B0000
0C000012
15000000
9461000C
A4630040
BC030000
10000005
15000000
9462000C
A8630040
DC02180C
9C21047C
A96E0000
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
03FFFFF0
9DC0FFFF
D7E117F4
D7E177F8
D7E14FFC
D7E10FF0
9C21FFF0
A9C30000
04000DFE
A8440000
BC0B0000
10000006
15000000
846B0038
BC230000
0C000044
15000000
98A2000C
A485FFFF
A4640008
BC030000
10000018
A4640010
84C20010
BC260000
0C000021
A4640280
A4640001
BC030000
10000026
A4840002
84620014
9C800000
E0601802
D4022008
D4021818
BC260000
0C000026
9D600000
9C210010
8521FFFC
8421FFF0
8441FFF4
44004800
85C1FFF8
BC230000
0C00003C
A4840004
BC240000
10000026
15000000
84C20010
A8850008
BC260000
DC02200C
13FFFFE4
A484FFFF
A4640280
BC030200
13FFFFE1
A4640001
A8820000
04000E2D
A86E0000
9482000C
03FFFFDA
84C20010
BC240000
10000003
15000000
84620014
D4021808
BC260000
13FFFFDE
9D600000
9862000C
A4830080
E4045800
13FFFFD9
A8630040
9D60FFFF
03FFFFD6
DC02180C
04000A7C
A86B0000
03FFFFBD
98A2000C
84820030
BC040000
1000000A
9C620040
E4041800
10000006
9C600000
04000AFC
A86E0000
98A2000C
9C600000
D4021830
84C20010
9C80FFDB
9C600000
E0A52003
D4021804
03FFFFCC
D4023000
9C600009
A8A50040
D40E1800
DC02280C
03FFFFB9
9D60FFFF
D7E117E8
18400001
D7E177EC
A8421D98
D7E197F0
85C20000
D7E1A7F4
850E0148
D7E1B7F8
D7E14FFC
D7E10FE4
BC280000
9C21FFE4
AAC30000
A8440000
AA850000
0C00003B
AA460000
84E80004
BD47001F
10000014
18600000
BC360000
10000025
9CA70001
9CE70002
D4082804
B8E70002
9D600000
E0E83800
D4071000
9C21001C
8521FFFC
8421FFE4
8441FFE8
85C1FFEC
8641FFF0
8681FFF4
44004800
86C1FFF8
A8630000
BC230000
0FFFFFF5
9D60FFFF
07FFE318
9C600190
BC0B0000
1000001F
A90B0000
846E0148
9C800000
D40B1800
D40B2004
D40E5948
D40B2188
D40B218C
BC360000
9CA00001
0FFFFFDF
A8E40000
B9670002
9C800001
BC360002
E0685800
E0843808
D403A088
84C80188
E0C62004
D4083188
13FFFFD4
D4039108
8468018C
E0832004
03FFFFD0
D408218C
9D0E014C
03FFFFC6
D40E4148
03FFFFD1
9D60FFFF
D7E117D8
18400001
D7E1F7F8
A8421D98
D7E197E0
87C20000
D7E1D7F0
D7E1E7F4
D7E14FFC
D7E10FD4
D7E177DC
D7E1A7E4
D7E1B7E8
D7E1C7EC
9C5E0148
9C21FFD0
1B800000
AB430000
AA440000
D4011000
AB9C0000
869E0148
BC340000
0C000043
86C10000
84540004
9DC2FFFF
BD6E0000
0C00002F
BC1C0000
9C420001
B8420002
0000000A
E0541000
84620100
E4039000
10000009
15000000
9DCEFFFF
BC2EFFFF
0C000022
9C42FFFC
BC120000
0FFFFFF7
15000000
84740004
9C63FFFF
E4237000
0C000041
84A20000
9C600000
D4021800
BC050000
13FFFFF1
9C600001
E0837008
84740188
E0641803
BC030000
0C00002C
87140004
48002800
15000000
84740004
E423C000
13FFFFD4
15000000
84760000
E423A000
13FFFFD0
9DCEFFFF
BC2EFFFF
13FFFFE2
9C42FFFC
BC1C0000
1000000F
15000000
84540004
BC220000
10000028
84540000
BC020000
10000025
A8740000
07FFE2A0
D4161000
86960000
BC340000
13FFFFC1
15000000
9C210030
8521FFFC
8421FFD4
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
8474018C
E0641803
BC230000
10000009
15000000
A87A0000
48002800
84820080
03FFFFD1
84740004
03FFFFC3
D4147004
48002800
84620080
03FFFFCB
84740004
AAD40000
03FFFFDF
AA820000
D7E117D8
84A30010
84440010
D7E1F7F8
D7E14FFC
D7E10FD4
D7E177DC
D7E197E0
D7E1A7E4
D7E1B7E8
D7E1C7EC
D7E1D7F0
D7E1E7F4
E5422800
9C21FFD4
1000007E
9FC00000
9C42FFFF
9F040014
BB820002
9E830014
AB440000
E1D8E000
E394E000
848E0000
AAC30000
9C840001
07FFF50B
847C0000
E40BF000
10000038
AA4B0000
A97E0000
A9140000
A8F80000
A89E0000
84670000
84C80000
A4A3FFFF
B8630050
E0A59306
E0639306
E0AB2800
A586FFFF
B9650050
E08C2000
A4A5FFFF
E16B1800
B8C60050
E0642802
A4ABFFFF
B8830090
E0C62802
A463FFFF
E0C62000
9CE70004
B8860010
E46E3800
B96B0050
E0641804
9D080004
D7E81FFC
13FFFFE6
B8860090
847C0000
BC230000
10000015
A8760000
9C7CFFFC
E4741800
1000000F
15000000
849CFFFC
BC240000
0C000008
9C63FFFC
0000000A
D4161010
84830000
BC040000
0C000005
9C63FFFC
E4741800
0FFFFFFB
9C42FFFF
D4161010
A8760000
0400140D
A89A0000
BD8B0000
10000032
A8F40000
9E520001
9CA00000
84C70000
84780000
A486FFFF
A503FFFF
E0A42800
B8630050
E0854002
B8C60050
B8A40090
A484FFFF
E0C61802
9F180004
E0C62800
9CE70004
B8660010
E46EC000
B8A60090
E0832004
13FFFFEE
D7E727FC
B8820002
E0942000
84640000
BC230000
10000017
ABD20000
9C64FFFC
E4741800
10000011
15000000
8484FFFC
BC240000
0C00000A
9C63FFFC
9C630004
0000000C
D4161010
84830000
BC040000
0C000006
15000000
9C63FFFC
E4741800
0FFFFFFA
9C42FFFF
D4161010
ABD20000
9C21002C
A97E0000
8521FFFC
8421FFD4
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
D7E117D8
D7E197E0
D7E1A7E4
D7E1B7E8
D7E1C7EC
D7E1F7F8
D7E14FFC
D7E10FD4
D7E177DC
D7E1D7F0
D7E1E7F4
85630040
9C21FF60
BC0B0000
D4013008
D4013818
D401401C
ABC30000
AAC40000
A8450000
870100A0
AA840000
1000000B
AA450000
84A30044
9C800001
D40B2804
E0A42808
A88B0000
04001132
D40B2808
9C600000
D41E1840
BD760000
0C000047
A9D60000
9CA00000
D4182800
18C07FF0
E06E3003
E4233000
0C000025
18800001
A9940000
A9A20000
A8841F78
84A40000
84C40004
E06C0004
E08D0004
04002694
AB820000
BC0B0000
0C00003B
8461001C
844100A4
BC020000
9C400001
19600001
D4031000
10000005
A96B1DD9
E04B1000
848100A4
D4041000
9C2100A0
8521FFFC
8421FFD4
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
BC220000
84E1001C
9C40270F
19600001
D4071000
1000000A
A96B1F71
1840000F
A842FFFF
E1CE1003
BC2E0000
10000005
844100A4
19600001
A96B1F68
844100A4
BC020000
13FFFFE2
15000000
904B0003
BC020000
0C000003
9C4B0008
9C4B0003
846100A4
03FFFFDA
D4031000
18807FFF
9C600001
A884FFFF
D4181800
E2962003
03FFFFB8
A9D40000
A8940000
A87E0000
A8A20000
9CC10070
9CE1006C
0400146C
BACE0054
BC160000
0C0001A8
D401582C
86C1006C
84A10070
E0B62800
BD85FBEF
100002A7
9C850412
9C60FC0E
E0632802
E0822048
E06E1808
E0632004
07FFF3D6
9DC5FFFF
1860FE10
9C800001
E16B1800
AB8C0000
D4012048
18600001
A9BC0000
A98B0000
A8631F80
84A30000
84C30004
E06C0004
E08D0004
07FFF0E1
15000000
18A00001
E06B0004
E08C0004
A8A51F88
84C50004
84A50000
07FFEEDE
15000000
18A00001
E06B0004
E08C0004
A8A51F90
84C50004
84A50000
04002341
15000000
D4015810
D4016014
0400277D
A86E0000
18A00001
E06B0004
E08C0004
A8A51F98
84C50004
84A50000
07FFEECA
15000000
84610010
84810014
E0AB0004
E0CC0004
0400232F
15000000
E06B0004
E08C0004
D4015810
D4016014
0400273F
15000000
18E00001
A8E71F78
84610010
84810014
84A70000
84C70004
040026BF
AB0B0000
BD8B0000
1000024F
9C600001
BC580016
10000014
D4011830
18A00001
B8780003
A8A52040
A8E20000
E0632800
A8D40000
84830004
84630000
E0A60004
E0C70004
04002632
15000000
BD4B0000
0C00024A
9CE00000
9CC00000
9F18FFFF
D4013030
E2D67002
9C600000
9F56FFFF
E57A1800
0C000230
D4011828
BD980000
10000225
9C800000
E35AC000
D401C040
D4012038
84610008
BC430009
1000013E
BDA30005
10000006
9C600001
84810008
9C600000
9C84FFFC
D4012008
84810008
BC040003
10000513
BD440003
0C0003B6
84C10008
BC060004
10000250
9CE00001
BC060005
0C0003B4
D4013834
84A10018
E0A5C000
9F850001
BD5C0000
0C000508
D401283C
BCBC000E
A8FC0000
10000003
9DC00001
9DC00000
E1C37003
9CC00000
BCA70017
D41E3044
1000000B
A8860000
9CA00001
9C600004
E0631800
A8850000
9CC30014
E4A63800
13FFFFFC
9CA50001
D41E2044
04001005
A87E0000
BC0E0000
D4015810
1000011C
D41E5840
BDB80000
D401A04C
100003AC
D4011050
A478000F
B9D80084
18E00001
B8630003
A8E72040
A48E0010
E0633800
BC040000
84830000
84A30004
D4012000
D4012804
10000379
A8940000
A9A20000
18400001
A9940000
A8422018
A5CE000F
84A20020
84C20024
E06C0004
E08D0004
07FFEB4E
9E400003
D4015820
D4016024
BC0E0000
10000014
18400001
85610000
85810004
A8422018
A48E0001
BC040000
E06B0004
E08C0004
10000006
B9CE0081
84A20000
84C20004
07FFEE2D
9E520001
BC2E0000
13FFFFF5
9C420008
D4015800
D4016004
84A10000
84C10004
84610020
84810024
07FFEB31
15000000
D4015800
D4016004
84410030
BC020000
1000000D
A8720000
18400001
84610000
84810004
A8421FA0
84A20000
84C20004
0400261D
15000000
BD8B0000
100004C3
A8720000
040026BA
18400001
E06B0004
E08C0004
84A10000
84C10004
07FFEE09
A8421FB0
84A20000
84C20004
E06B0004
E08C0004
0400226E
15000000
18A0FCC0
BC3C0000
A9CC0000
0C0002A4
E04B2800
D401C054
D401E044
84E10034
BC070000
10000379
84610044
9CA3FFFF
18E00001
B8A50003
A8E72040
18600001
E0A53800
84C10010
A8631FC0
9EC60001
84830004
84630000
84C50004
84A50000
07FFEAF8
15000000
A8EE0000
A8C20000
E06B0004
E08C0004
E0A60004
E0C70004
07FFEFDC
15000000
84610000
84810004
D4015820
D4016024
0400265C
15000000
A84B0000
A86B0000
04002682
9C420030
B8420018
84610000
84810004
E0AB0004
E0CC0004
07FFEFCB
B8420098
84E10010
D4015800
D4016004
D8071000
84610020
84810024
E0AB0004
E0CC0004
04002554
15000000
BD4B0000
10000067
18E00001
84A10000
84C10004
A8E71FA0
84670000
84870004
07FFEFB7
15000000
84610020
84810024
E0AB0004
E0CC0004
04002544
15000000
BD4B0000
1000022B
9C76FFFF
84410044
BDA20001
10000300
19C00001
84610010
A9CE1FA8
E0631000
868E0000
85CE0004
D401C060
D401D064
D401E068
AA560000
D4011844
D401A058
D401705C
AB830000
AB540000
00000012
AB0E0000
A8E71FA0
84670000
84870004
07FFEF95
15000000
84A10020
84C10024
E06B0004
E08C0004
0400259D
15000000
BD8B0000
10000208
E416E000
100002DD
15000000
A8EE0000
A8D40000
84610020
84810024
E0A60004
E0C70004
07FFED87
9ED60001
A8F80000
A8DA0000
84610000
84810004
E0A60004
E0C70004
D4015820
D4016024
07FFED7D
15000000
E06B0004
E08C0004
D4015800
D4016004
040025F8
15000000
A84B0000
A86B0000
0400261E
9C420030
B8420018
84610000
84810004
E0AB0004
E0CC0004
07FFEF67
B8420098
84A10020
84C10024
D8121000
D4015800
D4016004
E06B0004
E08C0004
0400256C
AA560000
BD8B0000
84A10000
84C10004
0FFFFFC1
18E00001
000000DD
87010054
18A0000F
18C03FF0
A8A5FFFF
9CE00000
E1742803
9DD6FC01
E16B3004
86C1006C
03FFFE64
D4013848
9C400000
A87E0000
D41E1044
A8820000
9C40FFFF
D401103C
04000EEF
9C400000
D4011018
9C400001
D4015810
D4011034
84410018
D41E5840
8781003C
D4011008
BDB8000E
84610070
10000003
9C400001
9C400000
A44200FF
BC020000
1000002C
BD830000
1000002A
15000000
18800001
B8780003
A8842040
BD5C0000
E0632000
84A30000
84C30004
D4012800
D4013004
1000010C
9C5CFFFF
84C10018
BD860000
0C000108
BC3C0000
100001ED
15000000
18400001
84610000
84810004
A8421FB8
84A20000
84C20004
07FFED1E
A9DC0000
A8F20000
A8D40000
E06B0004
E08C0004
E0A60004
E0C70004
040024A4
A85C0000
BD6B0000
0C000087
84A10010
84810018
86C10010
00000087
AF04FFFF
84410034
BC020000
0C0000C0
84410008
85C10038
86C10028
84410034
BDBA0000
1000000C
BDB60000
1000000A
E5BAB000
10000003
A87A0000
A8760000
84C10028
E2D61802
E0C61802
E35A1802
D4013028
84E10038
BDA70000
10000018
84610034
BC030000
10000394
BDAE0000
1000000E
A8820000
A87E0000
0400107A
A8AE0000
A87E0000
A88B0000
84A1002C
04000FE3
A84B0000
8481002C
A87E0000
04000EBB
D401582C
84810038
E0A47002
BC050000
0C0003BA
A87E0000
A87E0000
04000FC8
9C800001
84A10040
BDA50000
10000164
A9CB0000
A87E0000
04001062
A88B0000
84C10008
BDA60001
100003C9
A9CB0000
9CE00000
D4013800
846E0010
9C630004
B8630002
E06E1800
04000F43
84630000
9C600020
E1635802
E06BD000
A463001F
BC030000
100001EC
9C800020
E0841802
BDA40004
1000043C
84C10028
9C80001C
E0641802
E0C61800
E2D61800
D4013028
E35A1800
84610028
BDA30000
10000006
A87E0000
8481002C
0400109F
84A10028
D401582C
BDBA0000
10000006
A88E0000
A87E0000
04001098
A8BA0000
A9CB0000
84810030
BC040000
0C000284
84610008
BD430002
10000003
9C600001
9C600000
A46300FF
BC030000
10000169
BD5C0000
10000168
84E10034
BC3C0000
13FFFF89
9CA00005
A88E0000
A8DC0000
04000E79
A87E0000
8461002C
A88B0000
040010E1
A9CB0000
BD4B0000
0FFFFF7F
84810018
84A10010
9CC00031
9EC50001
D8053000
9F180001
A87E0000
04000E5C
A88E0000
BC220000
0C000006
A87E0000
A87E0000
04000E56
A8820000
A87E0000
8481002C
04000E52
9C580001
9CE00000
8461001C
D8163800
D4031000
844100A4
BC020000
100001C1
15000000
D402B000
03FFFD39
85610010
84A10028
E0C0C002
E0A5C002
9CE00000
D4012828
D4013038
03FFFDDA
D4013840
E340D002
D401D028
03FFFDD0
AB430000
0400250F
A8780000
84A10010
84C10014
E06B0004
E08C0004
040023AA
15000000
BC2B0000
0FFFFDAA
9C600001
03FFFDA8
9F18FFFF
03FFFDBB
D4013830
9C60FBEE
E0632802
03FFFD5E
E0621808
9C400001
D401E03C
D4011034
9C400000
D4011018
84410008
BD420001
0C00034A
9C5CFFFF
84610038
E5831000
0C000009
E1C31002
84810038
84A10040
E0622002
9DC00000
E0A51800
D4011038
D4012840
BD7C0000
0C000344
15000000
86C10028
A85C0000
84A10028
A87E0000
E0A51000
9C800001
D4012828
04000F1D
E35A1000
03FFFF2B
A84B0000
9CA00001
D4012834
84C10018
BDA60000
100002C6
BCA6000E
A8E60000
10000003
9DC00001
9DC00000
E1C37003
84610018
D401183C
03FFFDB4
AB830000
A9B20000
A9940000
84E10010
E06C0004
E08D0004
84A10000
84C10004
07FFE928
9EC70001
E06B0004
E08C0004
04002496
A9D40000
A86B0000
040024BD
AB4B0000
84A10000
84C10004
E06B0004
E08C0004
07FFEC0C
15000000
A9F20000
E0AB0004
E0CC0004
E06E0004
E08F0004
07FFEE00
15000000
9CBA0030
84C10010
A88B0000
BC1C0001
D8062800
A86C0000
10000050
A9640000
19C00001
AA630000
AA440000
A9CE1FA8
E0720004
E0930004
84AE0000
84CE0004
07FFEBF3
15000000
18E00001
D4015808
D401600C
A8E71F78
E06B0004
E08C0004
84A70000
84C70004
04002335
15000000
BC0B0000
13FFFF67
84610010
AA560000
00000013
E0431000
84AE0000
84CE0004
07FFEBDF
AA560000
18E00001
D4015808
D401600C
A8E71F78
E06B0004
E08C0004
84A70000
84C70004
04002321
15000000
BC0B0000
13FFFF54
A87E0000
84610008
8481000C
84A10000
84C10004
07FFE8DB
9ED60001
E06B0004
E08C0004
04002449
15000000
A86B0000
04002470
AB4B0000
84A10000
84C10004
E06B0004
E08C0004
07FFEBBF
15000000
84610008
8481000C
E0AB0004
E0CC0004
07FFEDB4
15000000
9CDA0030
A8AC0000
A88B0000
E4121000
D8123000
E0640004
E0850004
0FFFFFCF
A8AB0000
A9650000
A8EC0000
A84B0000
A8CB0000
A86C0000
E0A60004
E0C70004
E0830004
E0620004
04002010
15000000
84610000
84810004
D4015808
D401600C
E0AB0004
E0CC0004
040023A6
15000000
BD8B0000
1000000F
15000000
84610000
84810004
84A10008
84C1000C
040022E0
15000000
BC0B0000
0FFFFF13
A87E0000
A45A0001
BC020000
13FFFF0F
15000000
9056FFFF
D401C054
9C76FFFF
84A10010
00000008
A8830000
E4051800
1000022A
84410054
90440000
AAC30000
9C63FFFF
BC020039
13FFFFF9
9C84FFFF
9C420001
87010054
B8420018
B8420098
03FFFEF9
D8031000
84610008
9C800000
BD430001
0C00016F
D4012000
84A10040
BC050000
13FFFEA8
9D600001
03FFFE9F
846E0010
04002416
18400001
E06B0004
E08C0004
84A10000
84C10004
07FFEB65
A8421FB0
84A20000
84C20004
E06B0004
E08C0004
04001FCA
15000000
1860FCC0
A9CC0000
E04B1800
18A00001
84610000
84810004
A8A51FB8
84C50004
84A50000
07FFED4F
15000000
A8EE0000
A8C20000
D4015800
D4016004
E06B0004
E08C0004
E0A60004
E0C70004
040022D8
15000000
BD4B0000
100000C5
18C08000
A8EE0000
E0423000
84610000
84810004
A8C20000
E0A60004
E0C70004
04002347
15000000
BD8B0000
0C00008C
15000000
9DC00000
03FFFE27
A84E0000
84E10034
BC270000
1000015B
BDB60000
9E400000
8681002C
00000005
86C10010
04000D11
15000000
AA8B0000
A8740000
07FFFB15
A88E0000
E0769000
9D6B0030
9E520001
D8035800
E592E000
A87E0000
A8940000
9CA0000A
13FFFFF2
9CC00000
D4015818
E55C3000
0C000271
D401A02C
84610010
E2C3E000
9F800000
9CA00001
A87E0000
04000F01
8481002C
A88E0000
A86B0000
04000F60
D401582C
BD4B0000
0C000025
BC2B0000
90B6FFFF
9C76FFFF
84C10010
00000008
A8830000
E4061800
10000202
84A10010
90A40000
AAC30000
9C63FFFF
BC050039
13FFFFF9
9C84FFFF
9CA50001
D8032800
A87E0000
04000CD0
A88E0000
BC020000
13FFFE79
E07C1005
E0801802
E0641804
BD630000
13FFFE71
E060E002
E07C1804
BD630000
13FFFE6D
A87E0000
04000CC2
A89C0000
03FFFE6A
A87E0000
1000000B
9C76FFFF
84810018
A4640001
BC030000
10000005
15000000
03FFFFD7
90B6FFFF
AAC30000
9C76FFFF
90830000
BC040030
13FFFFFC
15000000
03FFFFDF
A87E0000
9C60001C
84E10028
E2D61800
E0E71800
E35A1800
03FFFE1B
D4013828
A8A20000
D4012020
D4012824
03FFFC93
9E400002
9CA00000
BC040002
13FFFE9D
D4012834
9C800000
A87E0000
D41E2044
04000C6A
9C400001
BDB8000E
D4015810
D41E5840
10000003
84610070
9C400000
A44200FF
BC020000
13FFFE6A
9F80FFFF
BD630000
0FFFFE67
9C400000
03FFFD81
D4011018
03FFFB7B
85610010
87010060
87410064
87810068
8681004C
03FFFD6E
86410050
E080C002
BC040000
10000157
A8A20000
A4A4000F
18600001
B8A50003
A8632040
A8E20000
A8D40000
B8440084
E0A51800
E0660004
E0870004
84C50004
84A50000
07FFEA9C
15000000
BC020000
D4015800
D4016004
13FFFC79
9E400002
19C00001
A9CE2018
A4820001
BC040000
E06B0004
E08C0004
10000006
B8420081
84AE0000
84CE0004
07FFEA8B
9E520001
BC220000
13FFFFF5
9DCE0008
D4015800
D4016004
03FFFC67
84410030
9DC00000
03FFFDF4
A84E0000
9E83FFFF
18800001
B8740003
A8842040
A8EE0000
A8C20000
E0432000
E0A60004
E0C70004
84620000
84820004
07FFEA74
15000000
84610000
84810004
D4015820
D4016024
040022EF
15000000
84A10010
A86B0000
A84B0000
04002314
9EC50001
84610000
84810004
E0AB0004
E0CC0004
07FFEC5E
9C420030
84C10044
84E10010
BC260001
D8071000
D4015800
D4016004
0C000025
84610010
84810044
A8560000
E2432000
84610000
84810004
18E00001
A8E71FA8
84A70000
84C70004
07FFEA50
9C420001
E06B0004
E08C0004
D4015800
D4016004
040022CB
15000000
A9CB0000
A86B0000
040022F1
9DCE0030
84610000
84810004
E0AB0004
E0CC0004
07FFEC3B
15000000
E4229000
E06B0004
E08C0004
13FFFFE7
DBE277FF
E2D6A000
D4015800
D4016004
18400001
84610020
84810024
A8421FC0
84A20000
84C20004
04001E9B
15000000
84A10000
84C10004
E06B0004
E08C0004
04002233
15000000
BD8B0000
0C000104
15000000
03FFFE9C
9056FFFF
8461002C
04000E71
A88E0000
BD6B0000
13FFFD7A
84610008
9CA0000A
A87E0000
8481002C
9CC00000
04000BFC
9F18FFFF
84A10034
BC050000
0C000027
D401582C
84A10008
BD450002
10000004
9C600001
84C10034
A8660000
A46300FF
BC030000
10000005
84E1003C
BDA70000
13FFFD6D
AB870000
03FFFED4
8781003C
E4322000
13FFFE93
84A10040
18C0000F
9CA00000
A8C6FFFF
E0743003
E4232800
13FFFE8B
D4012800
18E07FF0
E2943803
E4142800
13FFFE87
84A10040
84610028
9C800001
9C630001
9F5A0001
D4011828
03FFFE7F
D4012000
A87E0000
A8820000
9CC00000
04000BCE
9CA0000A
84C10008
A84B0000
BD460002
10000003
9C600001
9C600000
A46300FF
BC030000
10000006
15000000
84E1003C
BDA70000
13FFFD42
AB870000
8781003C
BDB60000
10000006
A8820000
A87E0000
04000DC2
A8B60000
A84B0000
84610000
BC030000
0C0000DD
AB420000
9F9CFFFF
86810010
A6520001
E394E000
D401C030
D401E028
AB0E0000
D4019020
85C1002C
A86E0000
07FFF9B0
A8980000
A86E0000
9CAB0030
A8820000
D4012818
04000E0E
D4015800
A87E0000
A8980000
A8BA0000
04000E29
AA4B0000
846B000C
BC230000
10000043
AACB0000
A86E0000
04000E02
A88B0000
AB8B0000
A87E0000
04000B84
A8960000
84C10008
E07C3004
BC230000
10000006
BD720000
84E10020
BC270000
0C0000FD
BD720000
0C0000C6
84E10008
E2523804
BC320000
10000006
BDBC0000
84610020
BC030000
100000FE
BDBC0000
0C0000DC
84C10018
84E10028
9E540001
D8143000
E4143800
100000E3
AAD20000
A88E0000
A87E0000
9CA0000A
04000B72
9CC00000
E422D000
0C000010
A9CB0000
A8820000
9CA0000A
9CC00000
A87E0000
04000B69
AA920000
A89A0000
A87E0000
9CA0000A
9CC00000
04000B63
A84B0000
03FFFFB8
AB4B0000
A8820000
A87E0000
9CA0000A
9CC00000
04000B5B
AA920000
A84B0000
03FFFFAF
AB4B0000
03FFFFC3
9F800001
9C800000
03FFFAF6
D4012034
BCBC000E
10000003
9DC00001
9DC00000
A5CE00FF
9C800000
E1CE1803
03FFFB07
D41E2044
9DC00001
D401703C
AB8E0000
03FFFFF9
D4017018
A87E0000
8481002C
04000CE9
84A10038
03FFFC7D
D401582C
9CA00030
84810010
9F020001
9C400031
D8042800
03FFFCD6
D8031000
A8940000
D4012000
D4012804
03FFFB32
9E400002
BC1C0000
13FFFDE2
15000000
8441003C
BDA20000
13FFFE9A
19C00001
A9CE1FA8
84610000
84810004
84AE0000
84CE0004
07FFE942
9C58FFFF
9C720001
D4011054
18400001
D4015800
D4016004
040021E6
A8421FB0
84610000
84810004
E0AB0004
E0CC0004
07FFE935
15000000
84A20000
84C20004
E06B0004
E08C0004
04001D9A
15000000
1860FCC0
8481003C
E04B1800
A9CC0000
03FFFB2F
D4012044
04000CB2
8481002C
03FFFC46
D401582C
84620000
84820004
84A10020
84C10024
07FFEB1A
15000000
84A10000
84C10004
E06B0004
E08C0004
040020A7
15000000
BD4B0000
10000005
8681004C
03FFFBD4
86410050
AAC20000
9C56FFFF
90620000
BC030030
13FFFFFC
87010054
03FFFC8E
A87E0000
BC120000
13FFFF09
18C0000F
9C600000
03FFFC37
D4011800
9CC00031
9F180001
03FFFE06
D8053000
84410048
BC020000
1000001A
15000000
9C430433
85C10038
03FFFCC2
86C10028
84410028
E2C2E002
03FFFCBE
9C400000
A87E0000
04000A98
84820004
84A20010
9C6B000C
9CA50002
9C82000C
B8A50002
04000936
AA8B0000
A87E0000
A8940000
04000CD4
9CA00001
03FFFF17
AB4B0000
8461006C
9C400036
85C10038
E0421802
03FFFCA8
86C10028
D401702C
84A10018
A9D80000
D4012808
87010030
8641002C
BD5C0000
0C000012
9CA00001
A87E0000
04000CC0
8481002C
A88E0000
A86B0000
04000D1F
AA4B0000
BD4B0000
0C00003D
BC2B0000
84A10018
BC050039
10000041
15000000
9CC50001
D4013008
AB820000
84410008
9ED40001
D8141000
D401902C
03FFFDC4
A85A0000
84610018
D401702C
BC230039
A9D80000
0C000023
87010030
84A10018
9C650001
AB820000
9ED40001
D8141800
03FFFDB7
A85A0000
D401702C
AB820000
A9D80000
A85A0000
03FFFD96
87010030
03FFFD91
9F800001
84610018
D401702C
BC030039
A9D80000
1000000E
87010030
BDB20000
13FFFFEC
84810000
03FFFFEA
9C640031
D401702C
84C10018
A9D80000
D4013008
87010030
03FFFFC1
8641002C
AB820000
A85A0000
9C800039
9ED40001
D8142000
03FFFD87
9CA00039
13FFFFCB
84810018
A4640001
BC030000
13FFFFC8
AB820000
03FFFFC0
84A10018
AB820000
D401902C
03FFFFF1
A85A0000
BC040004
13FFFBCB
9C80003C
03FFFDAA
E0641802
D7E117EC
9844000C
D7E1A7F8
AA830000
A462FFFF
D7E177F0
A9C40000
A4830008
D7E14FFC
D7E10FE8
D7E197F4
BC240000
10000044
9C21FFE8
A8420800
846E0004
BD430000
0C0000A3
DC0E100C
856E0028
BC0B0000
10000073
A442FFFF
9C600000
A4A21000
86540000
A4A5FFFF
E4051800
1000009E
D4141800
84AE0050
A4420004
BC020000
1000000A
A8740000
846E0030
844E0004
BC030000
10000004
E0A51002
844E003C
E0A51002
A8740000
848E001C
48005800
9CC00000
BC2BFFFF
0C000062
9C60F7FF
984E000C
848E0010
E0421803
D40E2000
A4621000
DC0E100C
9C400000
E4231000
10000079
D40E1004
848E0030
BC040000
1000004B
D4149000
9C4E0040
E4041000
10000004
15000000
04000247
A8740000
9C800000
D40E2030
9C210018
A9640000
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
864E0010
BC120000
10000036
A4630003
844E0000
BC230000
D40E9000
E0429002
10000003
9C600000
846E0014
BDA20000
0C000007
D40E1808
0000002B
9D600000
BD420000
0C000028
9D600000
A8B20000
A8C20000
856E0024
A8740000
48005800
848E001C
BD4B0000
E0425802
13FFFFF5
E2525800
944E000C
A8420040
9D60FFFF
DC0E100C
9C210018
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
84540000
BC220000
0C000046
AC620016
E0801802
E0641804
BD630000
10000007
AC42001D
E0601002
E0431004
BD820000
13FFFFE8
15000000
D4149000
9D600000
9C210018
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
84940000
AC44001D
E0602002
E0A01002
E0632004
E0451004
AC63FFFF
AC42FFFF
B863005F
B842005F
E0431004
BC220000
10000007
AC840016
E0402002
E0822004
BD640000
0C000022
15000000
984E000C
9C80F7FF
84AE0010
E0422003
D40E2800
A4821000
DC0E100C
9C400000
E4241000
0FFFFF8E
D40E1004
BC230000
0FFFFF8B
15000000
03FFFF89
D40E5850
846E003C
BD430000
13FFFF5D
9D600000
03FFFFD2
9C210018
A8740000
848E001C
48005800
9CC00001
BC2BFFFF
0FFFFFBA
A8AB0000
944E000C
03FFFF5D
856E0028
944E000C
A8420040
03FFFFAB
DC0E100C
D7E117F4
D7E177F8
D7E14FFC
D7E10FF0
BC030000
9C21FFF0
A8430000
10000006
A9C40000
84830038
BC240000
0C00000F
15000000
986E000C
BC030000
10000005
9D600000
A8620000
07FFFF26
A88E0000
9C210010
8521FFFC
8421FFF0
8441FFF4
44004800
85C1FFF8
0400011D
15000000
03FFFFF2
986E000C
D7E117F8
D7E14FFC
D7E10FF4
BC230000
9C21FFF4
0C00000C
A8430000
04000449
15000000
A8820000
07FFFFD8
A86B0000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
18400001
18800000
A8421D98
A8849790
04000406
84620000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E10FFC
9C21FFFC
9D600000
9C210004
44004800
8421FFFC
D7E10FFC
9C21FFFC
9D600000
9C210004
44004800
8421FFFC
18800000
D7E14FFC
D7E10FF8
A884EE80
040003EF
9C21FFF8
9C210008
8521FFFC
44004800
8421FFF8
18800000
D7E1A7E4
A88498A8
AA830000
D7E14FFC
D7E117D8
D7E177DC
D7E197E0
D7E1B7E8
D7E1C7EC
D7E1D7F0
D7E1E7F4
D7E1F7F8
D7E10FD4
9C400000
D414203C
9C6302EC
9C800003
85D40004
9CC00004
D41412E0
D41422E4
D4141AE8
9C21FFD4
9C6E005C
A8820000
D40E1000
D40E1004
D40E1008
DC0E300C
D40E1064
DC0E100E
D40E1010
D40E1014
D40E1018
9CA00008
1B800000
1B400000
1B000000
0400084A
1AC00000
AB9CD6D4
AB5AD754
AB18D7E4
AAD6D84C
86540008
9FC00001
9CC00009
D40EE020
D40ED024
D40EC028
D40EB02C
D40E701C
9C72005C
A8820000
D4121000
D4121004
D4121008
DC12300C
D4121064
DC12F00E
D4121010
D4121014
D4121018
04000831
9CA00008
9C600012
85D4000C
9CC00002
D412E020
D412D024
D412C028
D412B02C
D412901C
D40E1000
D40E1004
D40E1008
DC0E180C
D40E1064
D40E1010
D40E1014
D40E1018
DC0E300E
9C6E005C
A8820000
0400081C
9CA00008
D40EE020
D40ED024
D40EC028
D40EB02C
D40E701C
D414F038
9C21002C
8521FFFC
8421FFD4
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
D7E117F0
D7E177F4
9C44FFFF
9DC00068
D7E197F8
E1C27306
D7E14FFC
D7E10FEC
AA440000
9C21FFEC
04000486
9C8E0074
BC0B0000
10000009
A84B0000
9C6B000C
9C800000
D40B9004
D40B2000
D40B1808
040007F3
9CAE0068
9C210014
A9620000
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
D7E117F0
18400001
D7E177F4
A8421D98
D7E197F8
85C20000
D7E14FFC
844E0038
D7E10FEC
BC220000
9C21FFEC
10000004
AA430000
07FFFF6B
A86E0000
9DCE02E0
84AE0004
9CA5FFFF
BD850000
10000011
844E0008
9862000C
BC030000
10000013
9C820074
00000007
9CA5FFFF
98C4FF98
BC060000
1000000E
9C60FFFF
9CA5FFFF
9C44FFF4
BC25FFFF
13FFFFF9
9C840068
844E0000
BC220000
0C000021
15000000
03FFFFE8
A9C20000
9C60FFFF
9C800000
DC02180E
9C600001
9CA00008
DC02180C
9C600000
D4021864
D4021800
D4021808
D4021804
D4021810
D4021814
D4021818
040007B1
9C62005C
9C600000
A9620000
D4021830
D4021834
D4021844
D4021848
9C210014
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
A8720000
07FFFF9A
9C800004
BC0B0000
10000004
D40E5800
03FFFFC3
A9CB0000
9C40000C
03FFFFF0
D4121000
18600001
18800000
A8631D98
D7E14FFC
D7E10FF8
A884EE80
9C21FFF8
04000308
84630000
9C210008
8521FFFC
44004800
8421FFF8
84830038
D7E14FFC
D7E10FF8
BC240000
10000004
9C21FFF8
07FFFF13
15000000
9C210008
8521FFFC
44004800
8421FFF8
D7E10FFC
9C21FFFC
9C210004
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C210004
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C210004
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C210004
44004800
8421FFFC
D7E14FFC
D7E10FF8
04000315
9C21FFF8
18800000
A86B0000
040002A6
A8849878
9C210008
8521FFFC
44004800
8421FFF8
D7E14FFC
D7E10FF8
04000309
9C21FFF8
18800000
A86B0000
0400029A
A8849890
9C210008
8521FFFC
44004800
8421FFF8
D7E1A7F8
1A800001
D7E117EC
D7E177F0
D7E197F4
D7E14FFC
D7E10FE8
9C21FFE8
AA94476C
A8440000
040007A2
AA430000
84740008
85C30004
9C60FFFC
E1CE1803
9C60F000
E04E1002
9C420FEF
E0421803
E0421800
BD420FFF
0C000009
A8720000
04001893
9C800000
84740008
E0637000
E42B1800
0C00000D
A8720000
040007B7
A8720000
9C210018
9D600000
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
04001881
E0801002
BC2BFFFF
0C000015
18800001
E1CE1002
A8844FD4
84B40008
84640000
A9CE0001
E0431002
D4057004
A8720000
0400079F
D4041000
9C210018
9D600001
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
A8720000
04001868
9C800000
84740008
E04B1802
BDA2000F
13FFFFD7
18800001
A8420001
A8844764
D4031004
84840000
18400001
E16B2002
A8424FD4
03FFFFCE
D4025800
D7E177F8
D7E14FFC
D7E10FF0
D7E117F4
BC040000
9C21FFF0
1000004F
A9C30000
04000751
A8440000
8462FFFC
9C80FFFE
19000001
E0A32003
9CE2FFF8
A908476C
E0C72800
85680008
84860004
E42B3000
9D60FFFC
A4630001
0C000063
E0845803
BC230000
1000000E
D4062004
8442FFF8
18600001
E0E71002
E0A51000
A8634774
84470008
E4021800
10000070
15000000
8467000C
D402180C
D4031008
E0462000
84420004
A4420001
BC020000
0C000011
A8650001
E0A52000
18800001
84460008
A8844774
E4022000
10000081
A8850001
8486000C
A8650001
D402200C
D4041008
E0472800
D4071804
00000005
D4022800
E0472800
D4071804
D4022800
BC4501FF
1000001B
B8450049
B8A50043
9C800001
84680004
E0452800
B8A50082
B8420002
E0A42808
18800001
A884476C
E0A51804
E0422000
D4082804
84820008
D407100C
D4072008
D4023808
D404380C
04000730
A86E0000
9C210010
8521FFFC
8421FFF0
8441FFF4
44004800
85C1FFF8
BC420004
1000004A
BC420014
B8450046
9C620038
E0431800
19600001
B8420002
A96B476C
E0425800
84820008
E4241000
0C000044
15000000
84C40004
9C60FFFC
E0C61803
E4462800
0C000006
15000000
84840008
E4222000
13FFFFF8
15000000
84A4000C
D407280C
D4072008
D4053808
03FFFFDC
D404380C
BC230000
10000009
E0A42800
8442FFF8
E0E71002
E0A51000
84670008
8447000C
D403100C
D4021808
18400001
A8650001
A8424768
D4071804
84420000
E4651000
0FFFFFCA
D4083808
18400001
A86E0000
A8425004
07FFFF1F
84820000
03FFFFC3
15000000
E0462000
84420004
A4420001
BC020000
0C00000C
E0472800
8446000C
84660008
E0852000
D403100C
A8A40001
D4021808
E0472000
D4072804
03FFFFB3
D4022000
A8650001
D4071804
03FFFFAF
D4022800
10000015
BC420054
9C62005B
03FFFFB8
E0431800
B8430082
9C600001
84C80004
E0431008
A8A40000
E0423004
03FFFFC3
D4081004
D4083814
D4083810
E0672800
D407100C
D4071008
D4072004
03FFFF9A
D4032800
10000006
BC420154
B845004C
9C62006E
03FFFFA2
E0431800
10000006
BC420554
B845004F
9C620077
03FFFF9C
E0431800
10000006
15000000
B8450052
9C62007C
03FFFF96
E0431800
9C4000FC
03FFFF93
9C60007E
84C50008
D7E14FFC
D7E10FD4
D7E117D8
D7E177DC
D7E197E0
D7E1A7E4
D7E1B7E8
D7E1C7EC
D7E1D7F0
D7E1E7F4
D7E1F7F8
BC260000
0C00002C
9C21FFCC
94C4000C
ABC30000
A4660008
A8440000
BC030000
10000033
AA850000
84640010
BC230000
0C00002F
A6460002
A652FFFF
BC120000
10000037
85D40000
9EC00000
1B007FFF
AA560000
AB18FC00
BC120000
A8B60000
A87E0000
10000074
A8D20000
18807FFF
A884FC00
E4B22000
10000003
8482001C
A8D80000
85620024
48005800
15000000
BDAB0000
1000007F
E2D65800
84740008
E2525802
E1635802
BC2B0000
13FFFFEB
D4145808
9D600000
9C210034
8521FFFC
8421FFD4
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
A87E0000
07FFF390
A8820000
BC2B0000
10000120
15000000
94C2000C
A6460002
A652FFFF
BC120000
0FFFFFCD
85D40000
A6C60001
BC160000
10000060
AB920000
D4019000
AAD20000
BC160000
1000003A
9C600000
84810000
BC240000
0C0000B7
A87C0000
E4B2B000
10000003
AB120000
AB160000
84C20014
84620008
AB580000
E0661800
D4011804
84620000
84810004
E5582000
10000003
9C800001
9C800000
A48400FF
BC040000
1000000B
E5983000
84A20010
E4432800
10000003
9C800001
9C800000
A48400FF
BC040000
0C0000D0
E5983000
10000082
A89C0000
85620024
A87E0000
8482001C
48005800
A8BC0000
BD4B0000
0C00002C
AB4B0000
E252D002
BC320000
0C000082
A87E0000
84740008
E39CD000
E063D002
E2D6D002
BC230000
0FFFFFAA
D4141808
BC160000
0FFFFFCA
9C600000
878E0000
86CE0004
D4011800
03FFFFC2
9DCE0008
86CE0000
864E0004
03FFFF87
9DCE0008
18607FFF
A863FFFF
E4B21800
10000005
A8720000
18800001
A8841FC8
84640000
040018BB
A8980000
E0D85B06
A87E0000
85620024
8482001C
48005800
A8B60000
BD4B0000
10000021
15000000
9862000C
A8630040
9D60FFFF
03FFFF87
DC02180C
AA560000
BC120000
10000022
15000000
A4660200
BC030000
10000022
87820008
E492E000
10000053
AB1C0000
A4660480
BC230000
1000005D
15000000
84620000
A8960000
04000500
A8B80000
84620008
84820000
E383E002
E304C000
D402E008
D402C000
A9720000
84740008
E2D65800
E0635802
E2525802
BC030000
13FFFF65
D4141808
BC120000
0FFFFFE2
94C2000C
86CE0000
864E0004
03FFFFDB
9DCE0008
84620000
84820010
E4432000
10000006
E4B2E000
87020014
E472C000
13FFFFB9
E4B2E000
10000003
AB120000
AB1C0000
A8960000
040004DC
A8B80000
84620008
84820000
E063C002
E084C000
D4021808
BC030000
10000004
D4022000
03FFFFDB
A9780000
A87E0000
07FFFC77
A8820000
BC2B0000
13FFFFB6
15000000
03FFFFD3
A9780000
A8B80000
040004C7
E252D002
84620008
84820000
E063C002
E304C000
D4021808
BC320000
13FFFF83
D402C000
A87E0000
07FFFC64
A8820000
BC0B0000
0FFFFFA3
15000000
03FFFF7B
D4019000
AB920000
84620000
03FFFFB2
AB120000
9C80000A
04000404
A8B60000
BC0B0000
1000004E
9D6B0001
9C600001
E24BE002
03FFFF43
D4011800
84620014
84820010
E3031800
87420000
E0781800
E35A2002
BB03005F
9CFA0001
E0781800
E0E79000
BB030081
E4783800
10000004
A8B80000
AB070000
A8A70000
A4C60400
BC060000
10000028
A87E0000
04000185
A8850000
BC2B0000
0C000037
AB8B0000
A86B0000
84820010
04000435
A8BA0000
9462000C
9C80FB7F
E0632003
A8630080
DC02180C
E07CD000
E358D002
D402E010
D402C014
D4021800
AB920000
D402D008
03FFFF7D
AB120000
A89C0000
0400047B
84A10004
84A20000
84810004
A87E0000
E0A52000
A8820000
07FFFC1C
D4022800
BC0B0000
0FFFFF5B
87410004
03FFFF30
E252D002
04000A49
15000000
BC2B0000
13FFFFE5
AB8B0000
A87E0000
07FFFDD1
84820010
9862000C
9C80FF7F
E0632003
9C80000C
03FFFF4C
D41E2000
9C800001
9E560001
03FFFEF7
D4012000
03FFFECF
9D60FFFF
9C80000C
9862000C
03FFFF42
D41E2000
D7E1B7F4
9EC302E0
D7E14FFC
D7E10FE0
D7E117E4
D7E177E8
D7E197EC
D7E1A7F0
D7E1C7F8
BC160000
1000002A
9C21FFE0
AB040000
9E800000
85D60004
9DCEFFFF
BD8E0000
10000014
86560008
9C52000C
9E52000E
94A20000
BCA50001
9DCEFFFF
10000009
9C62FFF4
98920000
BC04FFFF
10000006
BC2EFFFF
4800C000
15000000
E2945804
BC2EFFFF
9C420068
13FFFFF2
9E520068
86D60000
BC360000
13FFFFE7
15000000
9C210020
A9740000
8521FFFC
8421FFE0
8441FFE4
85C1FFE8
8641FFEC
8681FFF0
86C1FFF4
44004800
8701FFF8
03FFFFF5
AA960000
D7E1B7F4
9EC302E0
D7E14FFC
D7E10FE0
D7E117E4
D7E177E8
D7E197EC
D7E1A7F0
D7E1C7F8
BC160000
10000029
9C21FFE0
AB040000
AA830000
9E400000
85D60004
9DCEFFFF
BD8E0000
10000012
84560008
9C42000C
94A20000
BCA50001
9DCEFFFF
10000009
9C82FFF4
98A20002
BC05FFFF
10000005
A8740000
4800C000
15000000
E2525804
BC2EFFFF
13FFFFF3
9C420068
86D60000
BC360000
13FFFFE9
15000000
9C210020
A9720000
8521FFFC
8421FFE0
8441FFE4
85C1FFE8
8641FFEC
8681FFF0
86C1FFF4
44004800
8701FFF8
03FFFFF5
AA560000
00001638
15000000
D7E14FFC
D7E10FF4
D7E117F8
BC250000
0C00000A
9C21FFF4
18800001
A8650000
A8841FCC
04000BBF
A8450000
BC0B0000
0C000009
18800001
19600001
A96B1D9C
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
A8620000
04000BB2
A8841D9C
BC0B0000
13FFFFF6
19600001
18800001
A8620000
04000BAB
A8841D9F
BC2B0000
0FFFFFEE
9D600000
03FFFFEF
9C21000C
D7E10FFC
9C21FFFC
19600001
9C210004
A96B4708
44004800
8421FFFC
18600001
D7E10FFC
A8634760
9C21FFFC
85630000
9C210004
44004800
8421FFFC
D7E10FFC
9C21FFFC
19600001
9C210004
A96B46E8
44004800
8421FFFC
D7E10FFC
9C21FFFC
9D600000
9C210004
44004800
8421FFFC
D7E10FFC
9C21FFFC
19600001
9C210004
A96B4728
44004800
8421FFFC
D7E14FFC
D7E117F4
D7E177F8
D7E10FF0
9C21FFF0
A9C30000
07FFFFB1
A8440000
A88E0000
A8A20000
07FFFFAF
A86B0000
9C210010
8521FFFC
8421FFF0
8441FFF4
44004800
85C1FFF8
D7E14FFC
D7E10FF8
07FFFFA3
9C21FFF8
9C210008
19600001
8521FFFC
A96B4728
44004800
8421FFF8
98A4000C
A4C5FFFF
D7E117EC
A4460002
D7E177F0
D7E14FFC
D7E10FE8
D7E197F4
D7E1A7F8
BC020000
9C21FFAC
0C00003B
A9C30000
A8440000
9884000E
BD840000
10000018
A4C60080
04001324
A8A10000
BD6B0000
0C000010
84810004
A8A08000
A484F000
AC642000
E4242800
E2401802
E2521804
AE52FFFF
0C000037
BA52005F
9462000C
A8630800
9E800400
0000000B
DC02180C
98A2000C
A4C5FFFF
A4C60080
BC060000
0C00002A
9E800400
A8A50800
9E400000
DC02280C
A86E0000
04000048
A8940000
BC2B0000
0C000039
18800000
9462000C
A8630080
A88498A8
BC120000
D40E203C
DC02180C
D4025800
D4025810
0C000025
D402A014
9C210054
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
9C440043
D4041000
D4041010
9C400001
D4041014
9C210054
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
03FFFFD8
9E800040
18800000
84620028
A884D7E4
E4232000
13FFFFC7
15000000
9462000C
9E800400
E063A004
D402A04C
03FFFFCF
DC02180C
9882000E
040012EC
A86E0000
BC0B0000
13FFFFD9
15000000
9462000C
A8630001
03FFFFD5
DC02180C
9862000C
A4830200
BC040000
0FFFFFD0
A8630002
9C820043
DC02180C
9C600001
D4022000
D4022010
03FFFFC9
D4021814
D7E177DC
9DC4000B
D7E197E0
D7E14FFC
D7E10FD4
D7E117D8
D7E1A7E4
D7E1B7E8
D7E1C7EC
D7E1D7F0
D7E1E7F4
D7E1F7F8
BCAE0016
9C21FFD0
10000035
AA430000
9C40FFF8
E1CE1003
B86E005F
BC230000
10000036
E4447000
10000003
9C400001
A8430000
A44200FF
BC020000
0C000030
9C40000C
040003B4
A8720000
BC4E01F7
1000002E
18800001
A884476C
E06E2000
8443000C
E4221800
0C00015F
B8AE0043
84820004
9CA0FFFC
8462000C
E0842803
84C20008
E0822000
D406180C
84A40004
D4033008
A8A50001
A8720000
040003C8
D4042804
9D620008
9C210030
8521FFFC
8421FFD4
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
BC440010
10000007
9C40000C
0400038B
9DC00010
03FFFFDA
18800001
9C40000C
9D600000
03FFFFEA
D4121000
B8AE0049
BC050000
1000008A
BC450004
100000BD
BC450014
B8AE0046
9CC50038
E0A63000
18E00001
B8A50002
A8E7476C
E0A53800
8445000C
E4051000
10000019
9D60FFFC
84620004
E0635803
E0837002
BD44000F
1000007A
BD640000
0C00000D
15000000
00000079
E0621800
9C80FFFC
84620004
E0632003
E0837002
BDA4000F
0C00006F
BD840000
0C00006F
15000000
8442000C
E4251000
13FFFFF5
15000000
9CA60001
1A800001
AA94476C
84540010
9D140008
E4224000
0C000107
9CC0FFFC
84620004
E0633003
E0837002
BDA4000F
0C0000F2
BD840000
D4144014
0C000066
D4144010
BC4301FF
10000090
B8830049
B8630043
9CE00001
84940004
E0C31800
B8630082
B8C60002
E0671808
18E00001
A8E7476C
E0632004
E0C63800
D4141804
84E60008
D402300C
D4023808
D4061008
D407100C
B8450082
9CC00001
E0C61008
E4461800
10000054
E0433003
BC220000
1000000F
E1652800
9C40FFFC
E0C63000
E0A51003
E0433003
BC220000
10000007
9CA50004
E0C63000
E0433003
BC020000
13FFFFFD
9CA50004
E1652800
18600001
B96B0002
A863476C
A9A50000
E16B1800
9D8B000C
9CECFFF4
844C0000
E4023800
10000019
9C80FFFC
84620004
E0632003
E0837002
BD44000F
100000CC
BD640000
0C00000D
E0821800
000000D2
84C2000C
9C80FFFC
84620004
E0632003
E0837002
BDA4000F
0C0000C1
BD840000
0C0000C7
15000000
8442000C
E4223800
13FFFFF5
15000000
9DAD0001
A44D0003
BC220000
13FFFFE1
9D8C0008
000000D5
A4650003
9CA0007E
03FFFF7C
9CC0003F
03FFFF99
9CC6FFFF
E0621800
84A2000C
84830004
84C20008
A8840001
D406280C
D4053008
D4032004
04000314
A8720000
03FFFF4D
9D620008
E0821800
A8720000
84A40004
A8A50001
0400030C
D4042804
03FFFF45
9D620008
84540008
9CA0FFFC
87020004
E3182803
E0787002
BDA3000F
10000003
9C800001
9C800000
A48400FF
BC240000
1000003A
E4987000
0C0000A2
9CA00001
A4A500FF
BC050000
0C000034
A88E0001
E1C27000
D4022004
A8630001
D4147008
D40E1804
040002F0
A8720000
03FFFF29
9D620008
0C000091
9CC5005B
BC450054
10000105
BC450154
B8AE004C
9CC5006E
03FFFF41
E0A63000
BC440004
0C00008B
BC440014
10000118
BC440054
9CC4005B
E0E63000
19600001
B8E70002
A96B476C
E0E75800
84870008
E4243800
0C0000FB
B8C60082
84C40004
9D60FFFC
E0C65803
E4833000
0C000006
15000000
84840008
E4272000
13FFFFF8
15000000
84E4000C
84740004
D402380C
D4022008
D4071008
03FFFF65
D404100C
1BC00001
18800001
ABDE4764
A8845004
847E0000
86C40000
BC23FFFF
0C0000EE
E2CEB000
9ED6100F
9CC0F000
E2D63003
A8720000
0400138B
A8960000
BC2BFFFF
0C000014
AB4B0000
19600001
E062C000
A96B476C
E443D000
E0825805
E0A02002
E0852004
9CA00001
B884005F
0C000079
D4012000
A4A500FF
BC050000
10000077
84810000
BC240000
0C000075
1B800001
84540008
9CE0FFFC
84A20004
E0A53803
E0657002
BDA3000F
10000003
9C800001
9C800000
A48400FF
BC240000
10000009
E44E2800
10000003
9CA00001
A8A40000
A4A500FF
BC050000
13FFFF98
A88E0001
0400028B
A8720000
03FFFEC4
9D600000
A86E0001
E1C27000
D4021804
A8A40001
D4147014
D4147010
E06E2000
D40E400C
D40E4008
D40E2804
D4032000
0400027C
A8720000
03FFFEB5
9D620008
03FFFF18
84740004
9C620008
84420014
E4031000
13FFFEEF
9CA50002
03FFFE9F
84820004
A8CE0001
8462000C
84A20008
D4023004
D405180C
E1C27000
03FFFFE5
D4032808
E0821800
84C2000C
84A40004
84E20008
A8A50001
A8720000
D4042804
D407300C
0400025F
D4063808
03FFFE98
9D620008
03FFFEB7
E0A63000
03FFFF60
A8A40000
B8830046
9CC40038
03FFFF79
E0E63000
856B0000
E40B1000
0C0000B6
15000000
A4650003
9C4BFFF8
BC230000
13FFFFF9
9CA5FFFF
84540004
AC66FFFF
E0431003
D4141004
E0C63000
E4A61000
10000003
9C600001
9C600000
A46300FF
BC030000
13FFFF37
E0603002
E0633004
BD630000
13FFFF33
E0623003
BC230000
13FFFEED
A8AD0000
E0C63000
E0623003
BC030000
13FFFFFD
9CA50004
03FFFEE7
E1652800
03FFFF89
9CA00000
1B800001
E423D000
AB9C4FD4
849C0000
E0962000
0C000066
D41C2000
84BE0000
BC25FFFF
0C000070
E07A1802
E0841800
D41C2000
A47A0007
BC030000
10000006
9CA01000
E35A1802
9CA01008
9F5A0008
E0A51802
E09AB000
A8720000
A4840FFF
E2C52002
040012E9
A8960000
BC0BFFFF
1000005B
9C600001
E06BD002
E0761800
A8630001
849C0000
84A10000
E0962000
D414D008
D41A1804
BC050000
10000011
D41C2000
BC58000F
0C000025
9CC0FFF8
84A20004
9C78FFF4
A4A50001
E0633003
9CE00005
E0A32804
E0C21800
D4022804
D4063804
BCA3000F
0C000047
D4063808
18400001
A8425000
84620000
E4A41800
10000003
18600001
D4022000
A8634FFC
84430000
E4441000
0C00001F
84540008
84A20004
9D60FFFC
D4032000
03FFFF4B
E0A55803
10000010
BC450554
B8AE004F
9CC50077
03FFFE3C
E0A63000
9C400001
03FFFF52
D41A1004
9CE00001
84740004
E0C73008
A8E40000
E0661804
03FFFF0E
D4141804
1000001B
15000000
B8AE0052
9CC5007C
03FFFE2C
E0A63000
03FFFF17
9ED60010
84A20004
9CE0FFFC
03FFFF2F
E0A53803
1000001F
BC440154
B883004C
9CC4006E
03FFFEE8
E0E63000
A4A30FFF
BC250000
13FFFF9A
15000000
E056C000
84740008
A8420001
03FFFFC6
D4031004
9CA000FC
03FFFE14
9CC0007E
03FFFFAA
9EC00000
18600001
A8634764
03FFFF92
D403D000
9C820008
18400001
A8720000
07FFFA2A
A8424FD4
03FFFFB6
84820000
10000006
BC440554
B883004F
9CC40077
03FFFEC9
E0E63000
10000005
B8830052
9CC4007C
03FFFEC4
E0E63000
9CE000FC
03FFFEC1
9CC0007E
03FFFF55
84540004
A4C30003
D7E10FF8
D7E117FC
BC060000
9C21FFF8
1000004C
A4C400FF
BC050000
1000004B
9D65FFFF
8CA30000
E4053000
0C00000C
9C630001
9C63FFFF
00000026
9C210008
1000001F
15000000
8CA30000
E4253000
0C00001F
9D6BFFFF
9C630001
A4A30003
BC250000
13FFFFF7
BC0B0000
BCAB0003
0C00001C
BC0B0000
10000011
15000000
8C830000
E4043000
10000011
9C830001
00000006
E1635800
8CA4FFFF
E4253000
0C00000B
15000000
E4245800
A8640000
13FFFFFA
9C840001
9D600000
9C210008
8421FFF8
44004800
8441FFFC
9C210008
A9630000
8421FFF8
44004800
8441FFFC
A48400FF
B8A40008
E0852004
B8A40010
E0A52004
84830000
1840FEFE
E0852005
A842FEFF
E0E41000
AC84FFFF
18408080
E0872003
A8428080
E0841003
BC240000
13FFFFD6
BC0B0000
9D6BFFFC
BC4B0003
13FFFFF1
9C630004
03FFFFD0
BC0B0000
03FFFFCB
A9650000
03FFFFDD
A9650000
D7E10FF8
D7E117FC
BCA5000F
1000004C
9C21FFF8
E0C32004
A4C60003
BC260000
1000003B
A8C30000
9EE5FFF0
9CC40004
BAF70044
9E630004
9E240008
B9770004
9DE30008
9DA4000C
9D6B0014
9D83000C
E1645800
A9040000
A8E30000
86A80000
9CC60010
D407A800
E4265800
86A6FFF0
9D080010
D413A800
9CE70010
86B10000
9E730010
D40FA800
9E310010
86AD0000
9DEF0010
D40CA800
9DAD0010
13FFFFF0
9D8C0010
9CF70001
A565000F
B8E70004
BCAB0003
E0C33800
10000027
E0843800
A9860000
A9040000
A8EB0000
85A80000
9CE7FFFC
D40C6800
BC470003
9D8C0004
13FFFFFB
9D080004
9CEBFFFC
9C40FFFC
A4A50003
E0E71003
BC250000
9CE70004
E0C63800
0C000009
E0843800
E0A62800
8C440000
9CC60001
DBE617FF
E4262800
13FFFFFC
9C840001
9C210008
A9630000
8421FFF8
44004800
8441FFFC
A8C30000
BC250000
13FFFFF2
15000000
03FFFFF8
9C210008
03FFFFFB
A8AB0000
D7E10FF8
D7E117FC
E4A32000
10000015
9C21FFF8
E0C42800
E4633000
10000012
BCA5000F
E0832800
BC250000
0C000008
E0A42802
9CC6FFFF
8C460000
9C84FFFF
E4242800
13FFFFFC
D8041000
9C210008
A9630000
8421FFF8
44004800
8441FFFC
BCA5000F
0C000012
E0C32004
A8C30000
BC050000
13FFFFF6
15000000
E0A62800
8C440000
9CC60001
DBE617FF
E4262800
13FFFFFC
9C840001
9C210008
A9630000
8421FFF8
44004800
8441FFFC
A4C60003
BC260000
13FFFFF2
A8C30000
9EE5FFF0
9CC40004
BAF70044
9E630004
9E240008
BAB70004
9DE30008
9DA4000C
9EB50014
9D83000C
E2A4A800
A9040000
A8E30000
85680000
9CC60010
D4075800
E426A800
8566FFF0
9D080010
D4135800
9CE70010
85710000
9E730010
D40F5800
9E310010
856D0000
9DEF0010
D40C5800
9DAD0010
13FFFFF0
9D8C0010
9CF70001
A5A5000F
B8E70004
BCAD0003
E0C33800
10000014
E0843800
A9860000
A9040000
A8ED0000
85680000
9CE7FFFC
D40C5800
BC470003
9D8C0004
13FFFFFB
9D080004
9CEDFFFC
9C40FFFC
A4A50003
E0E71003
9CE70004
E0C63800
03FFFFB7
E0843800
03FFFFB5
A8AD0000
A4C30003
D7E10FF8
D7E117FC
BC060000
10000054
9C21FFF8
BC250000
0C00004C
9CA5FFFF
B9A40018
A8E30000
A8C30000
00000005
B9AD0098
BC050000
10000044
A8AC0000
9CC60001
D8076800
A5060003
9D85FFFF
BC280000
13FFFFF8
9CE70001
BCA50003
10000030
BC050000
A4E400FF
BCA5000F
B9070008
E0E83804
B9070010
1000001B
E0E83804
9E25FFF0
9D060004
BA310044
9DE60008
9DA6000C
B9710004
A9860000
9D6B0014
E1665800
D40C3800
D4083800
9D080010
D40F3800
D40D3800
E4285800
9D8C0010
9DEF0010
13FFFFF8
9DAD0010
9E310001
A4A5000F
BA310004
BCA50003
1000000F
E0C68800
A9860000
A9050000
9D08FFFC
D40C3800
BC480003
13FFFFFD
9D8C0004
9CE5FFFC
9C40FFFC
A4A50003
E0E71003
9CE70004
E0C63800
BC050000
1000000A
15000000
B8840018
E0A62800
B8840098
D8062000
9CC60001
E4262800
13FFFFFD
15000000
9C210008
A9630000
8421FFF8
44004800
8441FFFC
03FFFFC0
A8C30000
D7E117F0
18400001
D7E177F4
D7E197F8
D7E14FFC
D7E10FEC
9C21FFEC
A8425010
040011A3
A9C30000
84620000
E4237000
0C00000C
AA4B0000
84820000
BC240000
13FFFFFE
18600001
A8AE0000
040011BF
A8635010
BC2B0000
13FFFFF8
15000000
18400001
A842500C
84620000
BC030000
0C000004
18600001
A8635014
D4039000
84620000
9C630001
D4021800
9C210014
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
18600001
D7E14FFC
A863500C
D7E10FF8
84830000
9C21FFF8
9C84FFFF
D4032000
84830000
BC240000
10000009
18600001
18A00001
A8635014
A8A55010
84630000
D4052000
0400117E
15000000
9C210008
8521FFFC
44004800
8421FFF8
84C3004C
D7E117F4
D7E177F8
D7E14FFC
D7E10FF0
BC260000
9C21FFF0
A8430000
0C000013
A9C40000
B8AE0002
E0A62800
85650000
BC0B0000
10000016
15000000
844B0000
D4051000
9C400000
D40B1010
D40B100C
9C210010
8521FFFC
8421FFF0
8441FFF4
44004800
85C1FFF8
9C800004
04000C0D
9CA00021
D402584C
BC2B0000
13FFFFEA
A8CB0000
03FFFFF3
9D600000
9C800001
A8620000
E0447008
9CA20005
04000C01
B8A50002
BC0B0000
13FFFFF7
15000000
D40B7004
03FFFFE4
D40B1008
D7E10FFC
BC040000
10000009
9C21FFFC
84A40004
84C3004C
B8650002
E0661800
84A30000
D4042800
D4032000
9C210004
44004800
8421FFFC
D7E117E8
D7E177EC
D7E197F0
D7E1A7F4
D7E14FFC
D7E10FE4
D7E1B7F8
A9C40000
84440010
9C21FFE4
AA430000
AA860000
9C840014
9D600000
84640000
9D6B0001
A4E3FFFF
B8630050
E0E72B06
E0632B06
E0C7A000
9C840004
B9060050
A4E6FFFF
E5425800
E1081800
B8C80010
BA880050
E0E63800
13FFFFF1
D7E43FFC
BC140000
1000000C
15000000
846E0008
E5821800
0C000012
A8720000
9C620005
9C420001
B8630002
E06E1800
D403A000
D40E1010
9C21001C
A96E0000
8521FFFC
8421FFE4
8441FFE8
85C1FFEC
8641FFF0
8681FFF4
44004800
86C1FFF8
848E0004
07FFFF8B
9C840001
84AE0010
9C8E000C
9CA50002
9C6B000C
B8A50002
07FFFE29
AACB0000
846E0004
8492004C
B8630002
E0641800
84830000
D40E2000
D4037000
03FFFFDF
A9D60000
D7E117E4
D7E177E8
D7E197EC
D7E1A7F0
D7E1B7F4
D7E14FFC
D7E10FE0
D7E1C7F8
AA430000
9C21FFE0
A8440000
9C660008
9C800009
AA860000
AAC50000
04001200
A9C70000
BDAB0001
10000038
9D000001
9C800000
E1084000
E54B4000
13FFFFFE
9C840001
07FFFF60
A8720000
9C600001
D40B7014
BDB60009
10000029
D40B1810
9F020009
E042B000
A9D80000
90CE0000
A8720000
A88B0000
9CA0000A
9CC6FFD0
07FFFF8F
9DCE0001
E42E1000
13FFFFF8
15000000
E058B000
9C42FFF8
E5B4B000
1000000D
E1D4B002
E1C27000
90C20000
A8720000
A88B0000
9CA0000A
9CC6FFD0
07FFFF7F
9C420001
E4227000
13FFFFF8
15000000
9C210020
8521FFFC
8421FFE0
8441FFE4
85C1FFE8
8641FFEC
8681FFF0
86C1FFF4
44004800
8701FFF8
9C42000A
03FFFFE7
9EC00009
03FFFFCF
9C800000
D7E117FC
1840FFFF
9C800000
E0A31003
D7E10FF8
E4252000
10000004
9C21FFF8
B8630010
9C800010
1840FF00
E0A31003
BC250000
10000004
1840F000
B8630008
9C840008
E0A31003
BC250000
10000004
1840C000
B8630004
9C840004
E0A31003
BC250000
10000005
BD830000
B8630002
9C840002
BD830000
10000010
15000000
18404000
E0631003
BC030000
0C000006
9D600020
9C210008
8421FFF8
44004800
8441FFFC
9C210008
9D640001
8421FFF8
44004800
8441FFFC
9C210008
A9640000
8421FFF8
44004800
8441FFFC
84830000
D7E10FFC
A4A40007
BC050000
1000000F
9C21FFFC
A4A40001
9D600000
E4255800
10000007
A4A40002
E4055800
0C00002D
9D600002
B8840042
D4032000
9C210004
44004800
8421FFFC
A4C4FFFF
BC260000
10000005
A4C400FF
B8840050
9CA00010
A4C400FF
BC260000
10000005
A4C4000F
B8840048
9CA50008
A4C4000F
BC260000
10000005
A4C40003
B8840044
9CA50004
A4C40003
BC260000
10000005
A4C40001
B8840042
9CA50002
A4C40001
BC260000
10000007
15000000
B8840041
BC040000
13FFFFDF
9D600020
9CA50001
9C210004
A9650000
D4032000
44004800
8421FFFC
B8840041
9C210004
9D600001
D4032000
44004800
8421FFFC
D7E14FFC
D7E117F8
D7E10FF4
A8440000
9C21FFF4
07FFFEB6
9C800001
9C800001
D40B1014
D40B2010
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E177EC
D7E1A7F4
85C40010
86850010
D7E197F0
D7E1B7F8
D7E14FFC
D7E10FE4
D7E117E8
E58EA000
9C21FFE4
AA440000
10000083
AAC50000
A8540000
AA8E0000
A9C20000
E0547000
84B20008
E5A22800
10000003
84920004
9C840001
07FFFE95
15000000
B9A20002
9DEB0014
E1AF6800
E48F6800
0C000007
A86F0000
9C800000
9C630004
E44D1800
13FFFFFE
D7E327FC
BA2E0002
9D960014
B9140002
E22C8800
9E720014
E48C8800
0C00004A
E1134000
872C0000
A779FFFF
BC1B0000
1000001F
BB390050
AAAF0000
AB330000
9CE00000
84790000
86F50000
A4C3FFFF
B8630050
E0C6DB06
E083DB06
A4B7FFFF
B8770050
E0A53000
9F390004
E0A53800
E0632000
B8E50050
A4A5FFFF
A8D50000
E0633800
9EB50004
B8830010
E448C800
B8E30050
E0A42804
13FFFFEB
D7F52FFC
D4063804
872C0000
BB390050
BC190000
10000021
AB6F0000
846F0000
AAB30000
AAEF0000
A8E30000
00000003
9CC00000
AB7D0000
84B50000
B8E70050
A4A5FFFF
A483FFFF
E0A5CB06
E0A53800
9EF70004
E0A53000
9EB50004
B8650010
9FBB0004
B8A50050
E0832004
E448A800
D7F727FC
9475FFFC
E063CB06
84FD0000
A487FFFF
E0632000
E0632800
13FFFFEA
B8C30050
D41B1804
9D8C0004
E4516000
13FFFFBA
9DEF0004
BD420000
0C000010
15000000
846DFFFC
BC230000
0C000008
9DADFFFC
0000000B
D40B1010
846D0000
BC030000
0C000006
15000000
9C42FFFF
BC020000
0FFFFFFA
9DADFFFC
D40B1010
9C21001C
8521FFFC
8421FFE4
8441FFE8
85C1FFEC
8641FFF0
8681FFF4
44004800
86C1FFF8
AA450000
03FFFF81
AAC40000
A4C50003
D7E117EC
D7E197F4
D7E1A7F8
D7E14FFC
D7E10FE8
D7E177F0
BC060000
9C21FFE8
A8450000
AA830000
0C000040
AA440000
B8420082
BC020000
10000029
15000000
85D40048
BC2E0000
0C000042
15000000
A4A20001
BC050000
0C00000F
15000000
B8420081
BC020000
1000001D
15000000
856E0000
BC2B0000
0C000022
A8AE0000
A9CB0000
A4A20001
BC050000
13FFFFF5
15000000
A8920000
A8AE0000
07FFFF46
A8740000
BC120000
1000001E
15000000
84920004
8474004C
B8840002
B8420081
E0832000
BC020000
84640000
D4121800
D4049000
0FFFFFE7
AA4B0000
9C210018
A9720000
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
A88E0000
07FFFF2C
A8740000
9CA00000
D40E5800
D40B2800
03FFFFDB
A9CB0000
03FFFFD0
AA4B0000
9CE6FFFF
18A00001
B8E70002
A8A51FE4
9CC00000
E0E72800
07FFFE07
84A70000
03FFFFBA
AA4B0000
A8740000
07FFFDC4
9C800001
9C600271
A9CB0000
D40B1814
9C600001
D40B1810
9C600000
D4145848
03FFFFB6
D40B1800
D7E1C7F8
BB050085
D7E1A7F0
86840010
D7E117E4
E298A000
84C40008
9C540001
D7E177E8
D7E197EC
D7E1B7F4
D7E14FFC
D7E10FE0
E5A23000
A9C40000
9C21FFE0
AAC50000
AA430000
10000006
84840004
E0C63000
E5423000
13FFFFFE
9C840001
07FFFDA1
A8720000
BDB80000
A90B0000
1000000C
9CEB0014
A8870000
9C600000
9C630001
9CA00000
E423C000
D4042800
13FFFFFC
9C840004
B8630002
E0E71800
84AE0010
A6D6001F
B8A50002
9CCE0014
BC160000
10000028
E0A62800
9D600020
9C800000
E16BB002
84660000
A9870000
E063B008
9CE70004
9CC60004
E0641804
E4453000
D7E71FFC
8466FFFC
13FFFFF7
E0835848
BC040000
10000003
D40C2004
9C540002
846E0004
8492004C
B8630002
9C42FFFF
A9680000
E0641800
D4081010
84430000
D40E1000
D4037000
9C210020
8521FFFC
8421FFE0
8441FFE4
85C1FFE8
8641FFEC
8681FFF0
86C1FFF4
44004800
8701FFF8
84660000
9CC60004
D4071800
E4453000
0FFFFFE8
9CE70004
84660000
9CC60004
D4071800
E4453000
13FFFFF6
9CE70004
03FFFFE1
846E0004
85630010
84A40010
D7E10FFC
E16B2802
BC2B0000
10000015
9C21FFFC
B8C50002
9C630014
9C840014
E0A33000
00000004
E0843000
0C000010
9D600000
9CA5FFFC
9C84FFFC
84E50000
84C40000
E4073000
13FFFFF9
E4832800
E4873000
10000003
9D60FFFF
9D600001
9C210004
44004800
8421FFFC
9C210004
44004800
8421FFFC
D7E177F0
A9C40000
D7E117EC
D7E197F4
D7E1A7F8
D7E14FFC
D7E10FE8
AA830000
9C21FFE8
A8850000
A86E0000
07FFFFD5
A8450000
BC2B0000
0C000058
AA4B0000
BD6B0000
0C000050
9E400000
A8740000
07FFFD22
848E0004
85EE0010
84C20010
BA2F0002
B8C60002
9C6E0014
9CA20014
D40B900C
E0853000
E2238800
9D8B0014
9CC00000
85030000
85A50000
A4E8FFFF
A44DFFFF
E0C73000
B9AD0050
E0E61002
B9080050
B8C70090
A4E7FFFF
E1086802
9CA50004
E0C83000
9DAC0004
B9060010
E4442800
9C630004
E0E83804
B8C60090
D40C3800
A84D0000
13FFFFEB
A98D0000
E4B11800
10000017
A8A30000
84830000
9D8C0004
A4E4FFFF
B8840050
E0C73000
9C630004
B8460090
A4E6FFFF
E4511800
E0C22000
B8460010
B8C60090
E0E23804
13FFFFF3
D7EC3FFC
AC45FFFF
9C60FFFC
E0428800
E0421803
9C420004
E04D1000
BC270000
10000007
9C42FFFC
9C42FFFC
84620000
BC030000
13FFFFFD
9DEFFFFF
D40B7810
9C210018
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
A86E0000
9E400001
A9C20000
03FFFFAF
A8430000
A8740000
07FFFCCF
A88B0000
9C600001
D40B9014
D40B1810
9C210018
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
D7E117FC
18407FF0
D7E10FF8
E0631003
1840FCC0
E0631000
BDA30000
1000000B
9C21FFF8
9C210008
9CA00000
A8C30000
A8E50000
8421FFF8
E1660004
E1870004
44004800
8441FFFC
E0601802
B8C30094
BD460013
0C000011
BD460032
9C600000
10000005
9C800001
9CA00033
E0C53002
E0843008
9C210008
A8A40000
A8C30000
A8E50000
8421FFF8
E1660004
E1870004
44004800
8441FFFC
18800008
9C210008
E0643088
9CA00000
8421FFF8
A8C30000
A8E50000
E1660004
E1870004
44004800
8441FFFC
D7E117E8
84430010
D7E177EC
B8420002
9DC30014
D7E197F0
E04E1000
D7E1A7F4
8642FFFC
D7E1B7F8
D7E14FFC
D7E10FE4
A8720000
9C21FFE4
07FFFD56
AA840000
9C600020
BD4B000A
E0635802
9EC2FFFC
1000001C
D4141800
9C60000B
18C03FF0
E0635802
E46EB000
E0B21848
9C800000
10000004
E0A53004
8482FFF8
E0841848
9D6B0015
E0525808
E0441004
9C21001C
A8E20000
A8C50000
8521FFFC
8421FFE4
E1660004
E1870004
8441FFE8
85C1FFEC
8641FFF0
8681FFF4
44004800
86C1FFF8
E46EB000
10000015
9CCBFFF5
BC060000
9CE2FFF8
10000014
8482FFF8
9C60002B
E0B23008
E1635802
E46E3800
E0645848
9CE00000
E0A51804
18603FF0
10000004
E0A51804
8442FFF4
E0E25848
E0443008
03FFFFDF
E0423804
BC260000
10000006
A8860000
18C03FF0
A8440000
03FFFFD8
E0B23004
E0B23008
9CE00000
18403FF0
A8870000
03FFFFF2
E0A51004
D7E117E4
D7E177E8
D7E197EC
D7E1A7F0
D7E1B7F4
D7E1C7F8
A9C40000
D7E14FFC
D7E10FE0
9C800001
9C21FFD8
AB050000
AAC60000
07FFFC31
AA870000
18607FFF
AA4B0000
A863FFFF
E04E1803
1860000F
B8420054
A863FFFF
BC220000
0C000004
E1CE1803
18600010
E1CE1804
BC180000
10000019
D4017004
A8610000
07FFFD25
D401C000
BC0B0000
0C000033
84610004
84810000
D4122014
D4121818
BC230000
10000003
9DC00002
9DC00001
BC020000
10000012
D4127010
9C42FBCD
9C600035
E0425800
E1635802
D4161000
00000017
D4145800
9C610004
07FFFD0E
9DC00001
84610004
D4127010
D4121814
BC020000
0FFFFFF2
9D6B0020
18603FFF
9D6BFBCE
A863FFFF
D4165800
E04E1800
B8420002
E0521000
84620014
07FFFCCB
B84E0005
E1625802
D4145800
9C210028
A9720000
8521FFFC
8421FFE0
8441FFE4
85C1FFE8
8641FFEC
8681FFF0
86C1FFF4
44004800
8701FFF8
9C800020
84A10000
E0845802
E0832008
E0635848
E0842804
D4011804
03FFFFCA
D4122014
D7E14FFC
D7E117EC
D7E177F0
D7E197F4
D7E1A7F8
D7E10FE8
9C21FFE0
AA440000
A8810000
07FFFF46
AA830000
A8720000
9C810004
A9CB0000
07FFFF41
A84C0000
84B40010
84920010
84610004
E0852002
84C10000
B8840005
E0C61802
E0662000
BDA30000
10000016
B8A30014
E0857000
A9C40000
A8A20000
A88E0000
A8CB0000
A8EC0000
E0640004
E0850004
E0A60004
E0C70004
07FFD725
15000000
9C210020
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
03FFFFEE
E16B2802
D7E177F8
D7E14FFC
D7E10FF0
D7E117F4
BD430017
9C21FFF0
0C00001E
A9C30000
18400001
A8421FD4
85620000
85820004
18800001
A84B0000
A86C0000
A8841FDC
84A40000
84C40004
E0830004
E0620004
07FFD9F6
9DCEFFFF
BC2E0000
13FFFFF6
18800001
A84B0000
9C210010
A8820000
A8AC0000
8521FFFC
8421FFF0
E1640004
E1850004
8441FFF4
44004800
85C1FFF8
18400001
B9C30003
A8422040
E1CE1000
844E0000
03FFFFF1
858E0004
9C84FFFF
84E50010
B9640085
B8E70002
9C850014
9D6B0001
E0E43800
B96B0002
D7E10FF8
D7E117FC
E4643800
9C21FFF8
10000015
E1635800
A8C30000
85040000
9C840004
D4064000
E4472000
13FFFFFC
9CC60004
E0872802
9C40FFFC
9C84FFEB
E0841003
9C840004
E0632000
E44B1800
0C000008
15000000
9C400000
9C630004
D7E317FC
E44B1800
13FFFFFC
15000000
9C210008
8421FFF8
44004800
8441FFFC
B8C40085
84A30010
D7E10FFC
E5653000
9C21FFFC
10000017
9C630014
B8850002
E0832000
E4632000
1000000F
9D600000
8564FFFC
BC2B0000
0C000008
9C84FFFC
0000001F
9C210004
84A40000
BC250000
1000001A
15000000
E4832000
13FFFFFB
9C84FFFC
9C210004
44004800
8421FFFC
E5453000
0C00000E
A4A4001F
BC250000
0C000012
B8860002
E0832000
84E40000
E0C72848
E0A62808
E4253800
13FFFFF2
9D600001
03FFFFE1
E4632000
B8860002
03FFFFDD
E0832000
9C210004
9D600001
44004800
8421FFFC
03FFFFD7
E0832000
D7E197E0
D7E1A7E4
D7E1C7EC
D7E14FFC
D7E10FD4
D7E117D8
D7E177DC
D7E1B7E8
D7E1D7F0
D7E1E7F4
D7E1F7F8
BC240000
9C21FFD4
AA440000
AB030000
0C0000B1
AA850000
07FFFAD6
9C54000B
84D2FFFC
9C60FFFC
BCA20016
9ED2FFF8
0C000052
E1C61803
9C800010
9CA00000
A8440000
E482A000
10000003
9C600001
9C600000
A46300FF
BC230000
100000A9
BC050000
0C0000A7
E56E2000
10000048
1B800001
E0767000
AB9C476C
84BC0008
E4051800
100000B5
9CE0FFFE
87830004
E0BC3803
E0A32800
84A50004
A4A50001
BC050000
0C000055
9CA0FFFC
E39C2803
E0BC7000
E5652000
1000008B
15000000
A4C60001
BC060000
0C000063
9CE0FFFC
8752FFF8
E356D002
84DA0004
E0C63803
E3853000
E57C2000
1000008A
9CAEFFFC
E3867000
E59C2000
10000058
A8940000
847A000C
849A0008
9CAEFFFC
D404180C
D4032008
BC450024
10000089
9C7A0008
BCA50013
1000000A
A8830000
84920000
BC45001B
D41A2008
84920004
100000E8
D41A200C
9C9A0010
9E520008
84B20000
AA830000
D4042800
A9DC0000
84720004
AADA0000
D4041804
84720008
D4041808
00000008
84DA0004
9C80FFF8
E0422003
A8820000
03FFFFB0
B8A2005F
AA920000
E06E1002
BCA3000F
0C000021
A4C60001
E0767000
E1C67004
D4167004
84430004
A8420001
D4031004
07FFFA98
A8780000
A9740000
9C21002C
8521FFFC
8421FFD4
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
A4C60001
BC060000
0C000015
9C60FFFC
8752FFF8
E356D002
84DA0004
03FFFFB7
E0C61803
E0961000
E0461004
A8A30001
D4161004
D4042804
E0441800
A8780000
84A20004
9C840008
A8A50001
07FFF2F2
D4022804
03FFFFDB
15000000
A8940000
07FFF675
A8780000
BC2B0000
0FFFFFD5
AA8B0000
84D2FFFC
9CA0FFFE
9C8BFFF8
E0662803
E0761800
E4241800
0C000090
9CAEFFFC
BC450024
1000007F
BCA50013
0C000068
BC45001B
A84B0000
A8720000
84830000
D4022000
84830004
D4022004
84630008
D4021808
A8920000
07FFF2D2
A8780000
03FFFFBB
15000000
07FFF656
A8850000
03FFFFBB
9C21002C
8483000C
84630008
AA920000
D403200C
D4041808
03FFFFA6
A9C50000
9C40000C
9D600000
03FFFFAF
D4181000
8483000C
84630008
D403200C
D4041808
847A000C
849A0008
BC450024
D404180C
D4032008
0FFFFF7B
9C7A0008
A8920000
07FFF949
AA830000
A9DC0000
84DA0004
03FFFF90
AADA0000
87C50004
9CE0FFFC
9C620010
E3DE3803
E3DE7000
E57E1800
1000003A
A4C60001
BC060000
0FFFFFB6
9CA0FFFC
8752FFF8
E356D002
84DA0004
E0C62803
E3DE3000
E5A3F000
0FFFFF55
9CAEFFFC
847A000C
849A0008
D404180C
D4032008
BC450024
10000060
9E9A0008
BCA50013
1000000A
A8740000
84720000
BC45001B
D41A1808
84720004
1000005C
D41A180C
9C7A0010
9E520008
84920000
D4032000
84920004
D4032004
84920008
D4032008
E07E1002
E09A1000
A8630001
D41C2008
D4041804
A8780000
849A0004
A4840001
E0422004
07FFF9FC
D41A1004
03FFFF65
A9740000
84520000
D40B1000
84520004
10000017
D40B1004
9C4B0008
03FFFF96
9C720008
E3DE1002
E2D61000
A87E0001
D41CB008
D4161804
A8780000
8492FFFC
A4840001
E0422004
07FFF9E7
D7F217FC
03FFFF50
A9720000
A86B0000
07FFF8F5
A8920000
03FFFF8B
A8920000
84520008
BC050024
D40B1008
8452000C
10000014
D40B100C
9C4B0010
03FFFF7B
9C720010
846BFFFC
9CE0FFFC
AA920000
E0633803
03FFFF2F
E1CE1800
84920008
BC050024
D41A2010
8492000C
1000000C
D41A2014
9C9A0018
03FFFF15
9E520010
84720010
9C4B0018
D40B1810
9C720018
84920014
03FFFF65
D40B2014
84B20010
9C9A0020
D41A2818
9E520018
84B2FFFC
03FFFF07
D41A281C
A8740000
07FFF8CA
A8920000
03FFFFB1
E07E1002
84720008
BC050024
D41A1810
8472000C
10000005
D41A1814
9C7A0018
03FFFFA1
9E520010
84920010
9C7A0020
D41A2018
9E520018
8492FFFC
03FFFF9A
D41A201C
E0A41804
D7E10FF8
D7E117FC
BC050000
9C21FFF8
0C000006
9D600002
9C210008
8421FFF8
44004800
8441FFFC
E0A02002
E0852004
AC84FFFF
B884005F
BC040000
10000008
18408000
E0A31000
E0C02802
E0A62804
BD650000
13FFFFF1
15000000
18407FFF
A842FFFF
E0631003
1840FFF0
E0A31000
18407FDF
A842FFFF
E4A51000
13FFFFE7
9D600004
1840000F
A842FFFF
E4A31000
13FFFFE2
9D600003
18407FF0
E0631005
E0A01802
E0651804
AC63FFFF
B863005F
03FFFFDA
E1641803
D7E117F8
A8440000
9884000E
D7E14FFC
D7E10FF4
04000876
9C21FFF4
BD8B0000
1000000A
9C80EFFF
84620050
E0635800
D4021850
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
9462000C
E0632003
DC02180C
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E10FFC
9C21FFFC
9D600000
9C210004
44004800
8421FFFC
98E4000C
D7E117EC
A8440000
A4870100
D7E177F0
D7E197F4
D7E1A7F8
D7E14FFC
D7E10FE8
BC040000
9C21FFE8
AA830000
AA450000
10000007
A9C60000
9882000E
9CA00000
04000837
9CC00002
98E2000C
9C60EFFF
9882000E
E0E71803
A8B20000
DC02380C
A8740000
040007B7
A8CE0000
9C210018
8521FFFC
8421FFE8
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
D7E117F8
A8440000
9884000E
D7E14FFC
D7E10FF4
0400081F
9C21FFF4
BC2BFFFF
0C00000A
9462000C
A8631000
D4025850
DC02180C
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
9C80EFFF
E0632003
DC02180C
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
9884000E
D7E14FFC
D7E10FF8
040007BC
9C21FFF8
9C210008
8521FFFC
44004800
8421FFF8
E1632004
D7E10FF8
A56B0003
D7E117FC
BC2B0000
10000024
9C21FFF8
84A30000
84C40000
E4253000
1000001F
1840FEFE
A842FEFF
E0C51000
ACA5FFFF
18408080
E0A62803
A8428080
E0A51003
BC250000
0C00000B
9C630004
9C63FFFC
0000002A
9C210008
18408080
A8428080
E0A51003
BC250000
10000027
9C630004
9C840004
1840FEFE
84C30000
85040000
A842FEFF
ACA6FFFF
E0E61000
E4064000
13FFFFF2
E0A72803
90A30000
BC050000
10000012
15000000
90C40000
E4262800
0C00000A
9C630001
9C63FFFF
0000000C
8C630000
90C40000
E4062800
0C000007
15000000
9C630001
90A30000
BC050000
0FFFFFF9
9C840001
8C630000
8D640000
E1635802
9C210008
8421FFF8
44004800
8441FFFC
9C210008
9D600000
8421FFF8
44004800
8441FFFC
D7E117DC
84440064
D7E1A7E8
A4422000
D7E1B7EC
D7E1C7F0
D7E14FFC
D7E10FD8
D7E177E0
D7E197E4
D7E1D7F4
D7E1E7F8
BC020000
9C21FFD8
AA840000
AAC30000
10000033
AB050000
84650008
87450000
BC230000
0C00002C
9F9A0004
865C0000
9DC00000
BA520042
E5527000
10000007
845A0000
0000001E
BA520002
E4327000
0C000019
15000000
84820000
A8760000
A8B40000
040005DF
9DCE0001
BC0BFFFF
0FFFFFF7
9C420004
9C400000
D4181008
D4181004
9C210028
8521FFFC
8421FFD8
8441FFDC
85C1FFE0
8641FFE4
8681FFE8
86C1FFEC
8701FFF0
8741FFF4
44004800
8781FFF8
84780008
BA520002
9F5A0008
9F9C0008
E0639002
BC230000
13FFFFD8
D4181808
03FFFFE9
9D600000
07FFF1CE
9C400000
03FFFFE7
D4181008
85650008
D7E14FFC
D7E10FF8
BC2B0000
0C000008
9C21FFF8
07FFFFB3
15000000
9C210008
8521FFFC
44004800
8421FFF8
9C210008
D4055804
8521FFFC
44004800
8421FFF8
D7E1A7E4
D7E14FFC
D7E10FD4
D7E117D8
D7E177DC
D7E197E0
D7E1B7E8
D7E1C7EC
D7E1D7F0
D7E1E7F4
D7E1F7F8
9C21FF2C
BC030000
D4011810
D4012004
D4013014
10000006
AA850000
84430038
BC220000
0C00026B
15000000
84410004
9862000C
A443FFFF
A4822000
BC240000
1000000A
9CA0DFFF
84410004
84820064
84E10004
A8432000
E0642803
DC07100C
D4071864
A442FFFF
A4620008
BC030000
1000022C
84810004
84640010
BC230000
0C000228
A442001A
BC22000A
0C000231
84E10004
9C400000
9E410068
D4011028
9C410067
9C600000
D4011000
D4019034
84A10000
D401183C
E0B22802
D4011838
A8520000
D401181C
D401282C
90740000
AC830025
A48400FF
BC040000
10000027
A9D40000
A46300FF
BC030000
0C000009
9DCE0001
9DCEFFFF
00000021
906E0000
BC230000
0C00000A
E2CEA002
9DCE0001
906E0000
AC830025
A48400FF
BC040000
0FFFFFF8
A46300FF
E2CEA002
BC160000
10000012
8481003C
84610038
E0962000
9C630001
D402A000
D402B004
D401203C
BD430007
0C00001F
D4011838
BC240000
10000354
84E1001C
D4012038
E0E7B000
A8520000
D401381C
906E0000
BC030000
10000137
9CC00000
9C600000
9DCE0001
D8011831
9F80FFFF
D4013008
ABC60000
908E0000
9E8E0001
9C64FFE0
BC430058
1000031A
18A00001
B8630002
A8A52108
E0632800
84630000
44001800
15000000
9C420008
84E1001C
E0E7B000
03FFFFE7
D401381C
ABDE0010
03FFFFEE
A9D40000
ABDE0010
A47E0010
BC030000
0C000291
84810014
A47E0040
BC030000
10000372
84610014
85C40000
9C630004
A5CEFFFF
D4011814
0000000C
9CA00001
ABDE0010
A4BE0010
BC050000
10000279
84810014
84A10014
9CA50004
D4012814
9CA00000
85C40000
9C800000
D401E020
D8012031
9EC00000
BD9C0000
10000003
9CE0FF7F
E3DE3803
E060E002
E063E004
BD830000
10000012
E0607002
E0637004
B863005F
BC030000
0C00000D
BC250000
100001CB
AB830000
A47E0001
BC030000
100001EA
15000000
9CA00030
8781002C
D8012867
00000018
9F010067
BC050001
100002E9
BC050002
10000056
AB120000
A46E0007
B9CE0043
9F18FFFF
9C630030
BC2E0000
13FFFFFB
D8181800
A49E0001
BC240000
0C000007
A8B80000
BC230030
0C000004
9C600030
9F18FFFF
DBE51FFF
E392C002
84810020
E57C2000
10000003
D401E00C
D401200C
BC160000
10000004
84A1000C
9CA50001
D401280C
A4FE0002
BC070000
10000005
D4013818
8461000C
9C630002
D401180C
A49E0084
BC040000
0C000046
D4012024
84A10008
84E1000C
E1C53802
BD4E0000
0C000040
BD4E0010
0C000348
8461003C
1AC00001
84C10038
AAD6227C
00000009
9F400010
9C860002
9C420008
A8C50000
9DCEFFF0
BD4E0010
0C000012
15000000
9CA60001
9C630010
D402B000
D402D004
D401183C
BD450007
0FFFFFF3
D4012838
BC230000
1000001C
A8C30000
9DCEFFF0
BD4E0010
9C800001
13FFFFF2
A8520000
E06E1800
D402B000
D4027004
D401183C
BD440007
10000172
D4012038
9C420008
0000001B
9CC40001
A46E000F
84810028
B9CE0044
E0641800
9F18FFFF
8C630000
BC2E0000
13FFFFF9
D8181800
03FFFFB4
E392C002
84610010
84810004
07FFFE85
9CA10034
BC2B0000
10000084
84C10038
8461003C
9C860001
03FFFFCE
A8520000
84810038
8461003C
9CC40001
90A10031
BC050000
1000000F
84A10018
9CA00001
9C810031
E0632800
D4022000
D4022804
D401183C
BD460007
10000130
D4013038
A8860000
9C420008
9CC60001
84A10018
BC050000
1000000F
84A10024
9C630002
9CE10032
9C800002
D4023800
D4022004
D401183C
BD460007
1000012D
D4013038
A8860000
9C420008
9CC60001
84A10024
BC250080
0C0000C8
84E10008
84E10020
E1C7E002
BDAE0000
10000028
1AC00001
BDAE0010
AAD6226C
0C00000B
9F400010
0000001A
E0637000
9CC40002
9C420008
A8850000
9DCEFFF0
BD4E0010
0C000012
15000000
9CA40001
9C630010
D402B000
D402D004
D401183C
BD450007
0FFFFFF3
D4012838
BC230000
10000029
9CC00001
9DCEFFF0
BD4E0010
A8830000
13FFFFF2
A8520000
E0637000
D402B000
D4027004
D401183C
BD460007
10000044
D4013038
9C420008
9CC60001
E063E000
D402C000
D402E004
D401183C
BD460007
0C000044
D4013038
BC230000
10000228
A45E0004
BC220000
10000108
D4011838
8441000C
84610008
E5621800
10000003
8481001C
A8430000
E0841000
D401201C
9C800000
A8520000
03FFFEA9
D4012038
84610010
84810004
07FFFE0F
9CA10034
BC2B0000
1000000E
84810038
8461003C
9CC40001
03FFFFC1
A8520000
8441003C
BC220000
0C000007
84A10004
84610010
84810004
07FFFE00
9CA10034
84A10004
9445000C
A4420040
BC220000
10000003
9D60FFFF
8561001C
9C2100D4
8521FFFC
8421FFD4
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
BC230000
10000217
9C400001
A87C0000
D4011038
D401C068
D401E06C
D401E03C
A8520000
9C420008
A49E0004
BC040000
1000002E
15000000
84810008
84A1000C
E1C42802
BDAE0000
10000028
15000000
BD4E0010
0C000275
15000000
1AC00001
84A10038
AAD6227C
00000009
9F000010
9CC50002
9C420008
A8A40000
9DCEFFF0
BD4E0010
0C000012
15000000
9C850001
9C630010
D402B000
D402C004
D401183C
BD440007
0FFFFFF3
D4012038
BC230000
10000024
9CC00001
9DCEFFF0
BD4E0010
A8A30000
13FFFFF2
A8520000
E0637000
D402B000
D4027004
D401183C
BDA60007
0C00018B
D4013038
8441000C
84E10008
E5623800
10000003
BC230000
A8470000
8461001C
E0631000
0FFFFF93
D401181C
84610010
84810004
07FFFDA4
9CA10034
BC2B0000
13FFFFA3
9C800000
A8520000
03FFFE34
D4012038
03FFFFA5
9D60FFFF
84610010
84810004
07FFFD98
9CA10034
BC2B0000
13FFFF97
84A10038
8461003C
9CC50001
03FFFFC6
A8520000
84A1000C
E1C72802
BDAE0000
13FFFF37
BDAE0010
1000022F
15000000
1AC00001
9F400010
00000009
AAD6226C
9CE40002
9C420008
A8850000
9DCEFFF0
BD4E0010
0C000012
15000000
9CA40001
9C630010
D402B000
D402D004
D401183C
BD450007
0FFFFFF3
D4012838
BC230000
10000014
9CE00001
9DCEFFF0
BD4E0010
A8830000
13FFFFF2
A8520000
E0637000
D402B000
D4027004
D401183C
BD470007
0C00014D
D4013838
BC230000
100001E8
9CC00001
A8830000
03FFFF0D
A8520000
84610010
84810004
07FFFD5E
9CA10034
BC2B0000
13FFFF5D
84810038
8461003C
9CE40001
03FFFFD6
A8520000
84610010
07FFE33D
84810004
BC0B0000
0FFFFFB5
84A10004
9445000C
A442001A
BC22000A
13FFFDD5
9C400000
84E10004
9847000E
BD820000
13FFFDD0
9C400000
84610010
A8870000
A8B40000
0400020D
84C10014
03FFFF4A
9C2100D4
BC230000
10000155
84410018
BC220000
0C000110
A8830000
9C600002
9CE10032
D401186C
D4013868
A8C50000
03FFFED7
A8520000
BC230000
10000153
9CC00001
A8830000
03FFFED4
A8520000
03FFFE56
AB120000
07FFEDDF
15000000
03FFFD96
84410004
BC230000
10000118
90410031
BC220000
0C00016F
A8830000
9C400001
9CA10031
A8C20000
D401106C
A8620000
D4012868
03FFFEAD
A8520000
84410008
8481000C
E1C22002
BD4E0000
13FFFF3D
A8520000
8441000C
84E10008
E5623800
0C00017F
15000000
8461001C
E0631000
03FFFEF5
D401181C
AB850000
03FFFE32
AB120000
84610014
84810014
84630000
9C840004
D4011808
BD630000
D4012014
13FFFDC9
A9D40000
E0601802
D4011808
ABDE0004
03FFFDC4
A9D40000
A9D40000
03FFFDC1
9CC0002B
9CE00000
A9140000
D4013808
9C64FFD0
84810008
9E940001
E0E42000
90880000
B8A70002
E0A72800
E0651800
D4011808
9C64FFD0
BCA30009
13FFFFF6
A9140000
03FFFDB2
9C64FFE0
ABDE0010
D8013031
A47E0010
BC030000
10000037
84810014
84A10014
9CA50004
D4012814
85C40000
BD8E0000
1000011F
9C80002D
92C10031
D401E020
03FFFDCF
9CA00001
18E00001
A47E0010
A8E71DB0
D8013031
D4013828
BC030000
10000077
84A10014
84610014
9C630004
D4011814
85C50000
A47E0001
BC030000
13FFFDBB
9CA00002
BC0E0000
13FFFDB8
9C600030
D8012033
D8011832
03FFFDB4
E3DE2804
84A10014
9CE00001
84650000
9CA50004
D8011840
9C600000
D401380C
D8011831
D4012814
AB870000
9F010040
9C800000
03FFFDE3
D4012020
A47E0010
D8013031
BC030000
0FFFFFCD
84810014
A47E0040
BC030000
10000112
84610014
84E10014
99C40002
9CE70004
03FFFFC8
D4013814
BC260000
13FFFD68
A9D40000
03FFFD66
9CC00020
ABDE0080
03FFFD63
A9D40000
A47E0040
BC030000
13FFFD87
84E10014
85C40000
9CE70004
A5CEFFFF
03FFFD87
D4013814
84E10014
9CA00001
9CE70004
D4013814
03FFFD81
85C40000
ABDE0001
03FFFD51
A9D40000
90940000
BC04002A
1000012F
9DD40001
9C64FFD0
AA8E0000
BCA30009
0C00000E
9CA00000
E0A52800
90940000
B8E50002
E0A53800
E0A32800
9C64FFD0
BCA30009
13FFFFF9
9E940001
BD650000
0C0000EA
15000000
03FFFD3C
AB850000
84E10014
18A00001
85C70000
A8A51DC1
9C600030
9C800078
9CE70004
D4012828
ABDE0002
D8011832
D8012033
D4013814
03FFFD59
9CA00002
ABDE0040
03FFFD29
A9D40000
18E00001
A47E0010
A8E71DC1
D8013031
D4013828
BC030000
0FFFFF8D
84A10014
A47E0040
BC030000
100000B0
84E10014
85C50000
84A10014
A5CEFFFF
9CA50004
03FFFF87
D4012814
A47E0010
BC030000
100000AA
D8013031
84A10014
84E1001C
84650000
9CA50004
D4033800
03FFFCD7
D4012814
84E10014
9C600000
87070000
D8011831
BC380000
0C0000CD
9F470004
BD9C0000
100000B3
A8780000
9C800000
07FFF35F
A8BC0000
BC0B0000
100000DA
9C800000
E38BC002
92C10031
D401D014
03FFFD57
D4012020
A8C50000
03FFFDD0
A8520000
BC230000
0FFFFF16
8441000C
84610010
84810004
07FFFC22
9CA10034
BC2B0000
13FFFE21
8461003C
03FFFE6E
8441000C
9C420008
9CC70001
03FFFDC4
A8870000
BC040000
13FFFE10
D8013031
9CE00001
9C600000
D401380C
D8012040
D8011831
AB870000
03FFFF5F
9F010040
84610010
84810004
07FFFC0A
9CA10034
BC2B0000
13FFFE09
84810038
8461003C
9CC40001
03FFFD8A
A8520000
BC4E0009
10000039
8781002C
9DCE0030
D8017067
03FFFD27
9F010067
84610010
84810004
07FFFBF8
9CA10034
BC2B0000
13FFFDF7
8461003C
03FFFE13
A8520000
84610010
84810004
07FFFBEF
9CA10034
BC2B0000
13FFFDEE
A8520000
03FFFCC3
84E1001C
84610010
84810004
07FFFBE6
9CA10034
BC2B0000
13FFFDE5
84810038
8461003C
9CC40001
03FFFD76
A8520000
84610010
84810004
07FFFBDB
9CA10034
BC2B0000
13FFFDDA
84810038
8461003C
9CC40001
03FFFD7B
A8520000
84610010
84810004
07FFFBD0
9CA10034
BC2B0000
13FFFDCF
84C10038
8461003C
9CC60001
03FFFD9F
A8520000
AB120000
A86E0000
9C80000A
07FFD001
9F18FFFF
9D6B0030
A86E0000
D8185800
07FFD806
9C80000A
BC2B0000
13FFFFF6
A9CB0000
03FFFCE5
E392C002
E1C07002
D8012031
D401E020
9EC0002D
03FFFCB0
9CA00001
84410018
BC220000
9CC00001
0FFFFD5A
A8520000
9C600002
9CA10032
D4121804
03FFFD4E
D4122800
84A10014
9CA50004
D4012814
9CA00001
03FFFC9C
85C40000
9CE70004
D4013814
03FFFEDB
85C50000
A47E0040
BC030000
1000000F
84E10014
84810014
84A1001C
84640000
9C840004
DC032800
03FFFC2B
D4012014
9C630004
D4011814
03FFFEB9
85C40000
03FFFE83
A8470000
8481001C
84670000
9CE70004
D4032000
03FFFC1F
D4013814
9CA0FFFF
03FFFC53
AB850000
07FFD8A9
D401D014
9CA00000
AB8B0000
92C10031
03FFFCAA
D4012820
84610010
84810004
07FFFB7B
9CA10034
BC2B0000
13FFFD7A
84810038
8461003C
9CC40001
03FFFD1F
A8520000
84810038
1AC00001
9C840001
03FFFCD3
AAD6227C
BCBC0006
10000003
A87C0000
9C600006
AB830000
AC63FFFF
1B000001
B863009F
D401D014
AB181DD2
E07C1803
03FFFEB3
D401180C
1AC00001
84C10038
AAD6227C
03FFFDA6
9CC60001
1AC00001
A8E60000
03FFFDEC
AAD6226C
92C10031
D401D014
03FFFC80
D4015820
84A10014
87850000
9CA50004
BD7C0000
13FFFC1A
D4012814
03FFFC18
9F80FFFF
D7E14FFC
D7E117F0
D7E177F4
D7E197F8
D7E10FEC
9C21FFEC
AA430000
A9C40000
07FFEF30
A8450000
A8920000
A8AE0000
A8C20000
07FFFB96
A86B0000
9C210014
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
94E4000C
D7E117F0
D7E177F4
A8440000
85C40064
9C80FFFD
D7E197F8
E0E72003
D7E14FFC
D7E10FEC
9C21FB84
9D000400
DC01380C
94E2000E
9D610068
85A2001C
85820024
DC01380E
A8810000
9CE00000
D4017064
AA430000
D401681C
D4016024
D4015800
D4015810
D4014008
D4014014
07FFFB71
D4013818
BD8B0000
10000008
A9CB0000
A8720000
07FFEA92
A8810000
BC0B0000
0C000012
15000000
9461000C
A4630040
BC030000
10000005
15000000
9462000C
A8630040
DC02180C
9C21047C
A96E0000
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
03FFFFF0
9DC0FFFF
E0842B06
D7E117F8
D7E14FFC
D7E10FF4
07FFEFC1
9C21FFF4
BC0B0000
1000000F
A84B0000
9C60FFFC
84ABFFFC
E0A51803
E0A51800
BC450024
1000001A
BCA50013
0C00000C
A86B0000
9C800000
D4032000
D4032004
D4032008
9C21000C
A9620000
8521FFFC
8421FFF4
44004800
8441FFF8
9C800000
BC45001B
D40B2000
0C000012
D40B2004
9C600000
BC050024
D40B1808
1000000F
D40B180C
03FFFFED
9C6B0010
A86B0000
07FFF313
9C800000
9C21000C
A9620000
8521FFFC
8421FFF4
44004800
8441FFF8
03FFFFE1
9C6B0008
9C6B0018
D40B2010
03FFFFDD
D40B2014
D7E177F4
D7E14FFC
D7E10FEC
D7E117F0
D7E197F8
BC240000
9C21FFEC
0C00000D
A9C30000
BC030000
10000006
A8440000
84830038
BC240000
0C00003F
15000000
9862000C
BC030000
0C00000A
A86E0000
9C210014
9D600000
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
07FFE960
A8820000
AA4B0000
8562002C
BC0B0000
10000007
A86E0000
48005800
8482001C
BD6B0000
0C00002B
15000000
9462000C
A4630080
BC030000
0C000028
A86E0000
84820030
BC040000
10000009
9C620040
E4041800
10000005
9C600000
07FFEBD2
A86E0000
9C600000
D4021830
84820044
BC040000
10000006
15000000
07FFEBCA
A86E0000
9C600000
D4021844
07FFEB47
15000000
9C600000
07FFEB49
DC02180C
9C210014
A9720000
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
07FFEB2E
15000000
03FFFFC2
9862000C
03FFFFD7
9E40FFFF
07FFEBB3
84820010
03FFFFD9
84820030
D7E14FFC
D7E117F8
D7E10FF4
9C21FFF4
07FFEE57
A8430000
A8820000
07FFFFA2
A86B0000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E117E8
D7E1A7F4
D7E1B7F8
D7E14FFC
D7E10FE4
D7E177EC
D7E197F0
9C21FFE0
AAC30000
AA840000
07FFEE70
A8450000
BC2B0001
0C00004D
9C74FFFF
A8760000
9C810003
A8B40000
040000FA
9CC2005C
BC2BFFFF
0C00002B
AA4B0000
BC2B0000
0C00002B
A9740000
90810003
0000000D
9DC00000
84620000
D8032000
84C20000
9CC60001
D4023000
9DCE0001
9C810003
E4B27000
10000019
E0647000
90830000
84C20008
9CC6FFFF
BD660000
13FFFFF2
D4023008
84620018
E5861800
1000001D
15000000
84620000
D8032000
84620000
8C830000
BC04000A
1000002C
9C630001
9DCE0001
D4021800
9C810003
E4B27000
0FFFFFEB
E0647000
00000005
A9740000
9462000C
A8630040
DC02180C
9C210020
8521FFFC
8421FFE4
8441FFE8
85C1FFEC
8641FFF0
8681FFF4
44004800
86C1FFF8
A8760000
A48400FF
04000045
A8A20000
AD6BFFFF
E0605802
E1635804
AD6BFFFF
B96B005F
BC2B0000
0FFFFFCD
9DCE0001
03FFFFEB
9D60FFFF
BC4300FE
13FFFFB5
A8760000
B8940018
AA4B0000
B8840098
03FFFFBB
D8012003
03FFFFEC
A8760000
98C5000C
A4E62000
D7E14FFC
D7E10FF8
BC270000
10000007
9C21FFF8
84E50064
A8C62000
A8E72000
DC05300C
D4053864
07FFFF90
15000000
9C210008
8521FFFC
44004800
8421FFF8
D7E117F0
D7E177F4
D7E197F8
D7E14FFC
D7E10FEC
9C21FFEC
AA430000
07FFEDD0
A9C40000
BC0B0000
10000008
A84B0000
846B0038
BC230000
10000005
A8620000
07FFEA90
A86B0000
A8620000
A8920000
07FFFFDA
A8AE0000
9C210014
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
D7E117F0
D7E177F4
D7E197F8
D7E14FFC
D7E10FEC
BC030000
9C21FFEC
AA430000
A9C40000
10000006
A8450000
84830038
BC240000
0C000056
15000000
98E2000C
A4C7FFFF
84A20018
A4660008
BC030000
10000045
D4022808
84A20010
BC250000
0C000042
A8720000
A4C62000
BC260000
0C000022
A5CE00FF
84620000
84820014
E0A32802
E5652000
10000027
15000000
9CA50001
84820008
9CC30001
9C84FFFF
D4023000
D4022008
D8037000
84620014
E4032800
10000024
BC2E000A
10000008
A96E0000
9462000C
A4630001
BC030000
0C00001E
A8720000
A96E0000
9C210014
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
84620064
9C80DFFF
A8E72000
E0632003
84820014
D4021864
84620000
E0A32802
E5652000
0FFFFFDD
DC02380C
A8720000
07FFE902
A8820000
BC2B0000
1000000A
9CA00001
03FFFFD6
84620000
A8720000
07FFE8FA
A8820000
BC2B0000
0FFFFFE1
15000000
03FFFFE0
9D60FFFF
A8720000
07FFDF5C
A8820000
BC0B0000
0FFFFFDA
9D60FFFF
98E2000C
84A20010
03FFFFB9
A4C7FFFF
07FFEA20
15000000
03FFFFAB
98E2000C
D7E14FFC
D7E117F4
D7E177F8
D7E10FF0
9C21FFF0
A9C30000
07FFED4D
A8440000
A88E0000
A8A20000
07FFFF8F
A86B0000
9C210010
8521FFFC
8421FFF0
8441FFF4
44004800
85C1FFF8
D7E117E8
D7E177EC
D7E197F0
D7E1A7F4
D7E14FFC
D7E10FE4
D7E1B7F8
A9C30000
BC240000
18600001
9C21FFD8
A8440000
A8634B74
AA850000
0C000019
AA460000
07FFED57
86C30000
A86E0000
A8820000
A8B40000
A8CB0000
4800B000
A8F20000
BC2BFFFF
10000005
9C400000
D4121000
9C40008A
D40E1000
9C210028
8521FFFC
8421FFE4
8441FFE8
85C1FFEC
8641FFF0
8681FFF4
44004800
86C1FFF8
07FFED40
86830000
A86E0000
A8810000
A8A20000
A8CB0000
4800A000
A8F20000
03FFFFEA
BC2BFFFF
D7E117E8
D7E177EC
D7E197F0
D7E1A7F4
D7E14FFC
D7E10FE4
D7E1B7F8
9C21FFD8
A8430000
AA840000
07FFED06
AA450000
18600001
BC220000
A9CB0000
0C000019
A8634B74
07FFED25
86C30000
A86E0000
A8820000
A8B40000
A8CB0000
4800B000
A8F20000
BC2BFFFF
10000005
9C400000
D4121000
9C40008A
D40E1000
9C210028
8521FFFC
8421FFE4
8441FFE8
85C1FFEC
8641FFF0
8681FFF4
44004800
86C1FFF8
07FFED0E
86830000
A86E0000
A8810000
A8A20000
A8CB0000
4800A000
A8F20000
03FFFFEA
BC2BFFFF
D7E10FFC
BC040000
1000000A
9C21FFFC
BCA500FF
0C00000B
9D60FFFF
D8042800
9D600001
9C210004
44004800
8421FFFC
9C210004
A9640000
44004800
8421FFFC
9C80008A
03FFFFF8
D4032000
D7E117E8
18400001
D7E14FFC
D7E177EC
D7E197F0
D7E1A7F4
D7E1B7F8
D7E10FE4
A8424B74
9C21FFE4
A9C60000
AAC30000
AA840000
AA450000
07FFECE3
84420000
A8760000
A8940000
A8B20000
A8EE0000
48001000
A8CB0000
9C21001C
8521FFFC
8421FFE4
8441FFE8
85C1FFEC
8641FFF0
8681FFF4
44004800
86C1FFF8
D7E117F0
D7E177F4
D7E197F8
D7E14FFC
D7E10FEC
BC260000
9C21FFEC
AA460000
A8450000
10000009
E1C53000
00000014
9C210014
0400010A
9C420001
E4227000
0C00000E
15000000
90620000
BC23000A
13FFFFF9
15000000
9C60000D
04000100
9C420001
040000FE
9062FFFF
E4227000
13FFFFF6
15000000
9C210014
A9720000
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
D7E14FFC
D7E10FF8
040003F9
9C21FFF8
15000000
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E14FFC
D7E10FF8
040003EA
9C21FFF8
9C600058
D40B1800
9C210008
9D60FFFF
8521FFFC
44004800
8421FFF8
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800058
9C210004
9D600000
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E14FFC
D7E10FF8
040003AF
9C21FFF8
9C600058
D40B1800
9C210008
9D60FFFF
8521FFFC
44004800
8421FFF8
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800058
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800005
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C800005
9C210004
9D60FFFF
D4032000
44004800
8421FFFC
18600001
D7E10FFC
A8630710
9C21FFFC
84630000
9C630002
8C630000
9C210004
44004800
8421FFFC
D7E117F4
18400001
D7E177F8
A8420710
D7E14FFC
85C20000
D7E10FF0
BC0E0000
1000002C
9C21FFF0
18600001
18A00001
A8630714
9CC00000
84830000
18600001
A8A55018
A863070C
B8840004
84630000
D4053000
07FFD43D
9DCE0003
9C60FF80
A48B00FF
D80E1800
A56BFFFF
84620000
9CC0FFC3
D8032000
B86B0048
84820000
9D600000
9C840001
D8041800
9C800003
84620000
9C630003
D8032000
84620000
9C630002
D8033000
9C600000
84420000
9C420001
D8021800
9C210010
8521FFFC
8421FFF0
8441FFF4
44004800
85C1FFF8
03FFFFFA
9D60FFFF
18800001
B8630018
A8840710
D7E10FFC
84C40000
B8630098
9C21FFFC
9CA60005
8C850000
A4840020
BC040000
13FFFFFD
15000000
A46300FF
D8061800
9C210004
44004800
8421FFFC
D7E117F8
18400001
D7E14FFC
A8420710
D7E10FF4
84820000
18400001
9C840001
A8425018
9C21FFF4
D4021800
9C400001
9CA00000
D8041000
18400001
18800000
A8420718
A884F940
040000DF
84620000
04000133
84620000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
18800001
A8840710
84840000
E4040000
10000004
15000000
03FFFFCD
15000000
44004800
15000004
B4600001
A4830004
E4040000
10000021
15000000
B4C00011
9CA0FFFF
ACA50010
E0A62803
C0002811
B4600006
A4830080
B8E40047
A9000010
E1C83808
A4830078
B8E40043
A9000001
E1A83808
9CC00000
E0AE3808
C0803002
E4262800
13FFFFFE
E0C67000
B4C00011
A8C60010
C0003011
15000000
15000000
15000000
15000000
15000000
15000000
15000000
15000000
B4600001
A4830002
E4040000
10000019
15000000
B4C00011
9CA0FFFF
ACA50008
E0A62803
C0002811
B4600005
A4830080
B8E40047
A9000010
E1C83808
A4830078
B8E40043
A9000001
E1A83808
9CC00000
E0AE3808
C0603003
E4262800
13FFFFFE
E0C67000
B4C00011
A8C60008
C0003011
44004800
15000000
B5A00011
A9AD0010
C0006811
15000000
15000000
15000000
15000000
15000000
44004800
15000000
B5A00011
9D80FFFF
AD8C0010
E18D6003
C0006011
44004800
15000000
44004800
C0801802
B5A00011
A9AD0008
C0006811
15000000
15000000
15000000
15000000
15000000
44004800
15000000
B5A00011
9D80FFFF
AD8C0008
E18D6003
C0006011
44004800
15000000
44004800
C0601803
D4011008
D4012814
D4013018
D401381C
D4014020
D4014824
D4015028
D401582C
D4016030
D4016834
D4017038
D401783C
D4018040
D4018844
D4019048
D401984C
D401A050
D401A854
D401B058
D401B85C
D401C060
D401C864
D401D068
D401D86C
D401E070
D401E874
D401F078
D401F87C
B5C00020
D4017080
B5C00040
D4017084
1A800001
AA944B80
86940000
1AA00001
AAB5512C
D415A000
A5A3FF00
B9AD0046
9DADFFF8
19C00001
A9CE5148
E1CE6800
85AE0000
E42D0000
0C000034
15000000
48006800
E0642004
1A800001
AA945130
86940000
1AA00001
AAB5512C
D415A000
18400001
A8425134
84620000
9C63FFFF
D4021800
84410080
C0001020
84410084
C0001040
84410008
8461000C
84810010
84A10014
84C10018
84E1001C
85010020
85210024
85410028
8561002C
85810030
85A10034
85C10038
85E1003C
86010040
86210044
86410048
8661004C
86810050
86A10054
86C10058
86E1005C
87010060
87210064
87410068
8761006C
87810070
87A10074
87C10078
87E1007C
84210004
24000000
15000000
07FFD388
E0642004
D7E117FC
18400001
B8630002
A842501C
D7E10FF8
E0C31000
18400001
9C21FFF8
A842509C
D4062000
E0631000
D4032800
9C210008
8421FFF8
44004800
8441FFFC
D7E10FFC
9C800011
9C21FFFC
B4640000
A8630004
C0041800
9C210004
44004800
8421FFFC
D7E10FF8
D7E117FC
9C600011
9C21FFF8
B5630000
9C40FFFB
E08B1003
C0032000
9C210008
B96B0042
8421FFF8
A56B0001
44004800
8441FFFC
D7E10FF8
D7E117FC
9C800011
9C21FFF8
B4840000
9C40FFFB
BC230000
E0841003
10000003
9CA00004
A8A30000
E0652004
9C800011
C0041800
9C210008
8421FFF8
44004800
8441FFFC
9C21FFFC
D4014800
B6804802
1A000001
AA10501C
1A400001
AA52509C
E094000F
E4240000
0C000010
15000000
9EC4FFFF
B8D60002
E1C68000
E1A69000
85CE0000
E42E0000
0C000004
15000000
48007000
846D0000
A8C00001
E0C6B008
03FFFFF0
E2943005
85210000
C120A002
44004800
9C210004
9C21FFFC
D4012000
A8800001
E0841808
B4604800
E0632004
C1201800
84810000
44004800
9C210004
9C21FFFC
D4012000
A8800001
E0841808
AC84FFFF
B4604800
E0632003
C1201800
84810000
44004800
9C210004
D7E14FFC
D7E117E4
D7E197EC
D7E1A7F0
D7E1B7F4
D7E1C7F8
D7E10FE0
D7E177E8
9C21FFE0
AA840000
07FFFFA4
18400001
04000170
AACB0000
18600001
A8424B7C
A863511C
9C800000
84A20000
AB0B0000
040000BF
AA430000
84520000
18600001
A8820000
A863511C
040000B9
E0B41000
E42B1000
13FFFFF9
A9CB0000
0400016B
A8780000
07FFFF9B
A8760000
9C210020
A96E0000
8521FFFC
8421FFE0
8441FFE4
85C1FFE8
8641FFEC
8681FFF0
86C1FFF4
44004800
8701FFF8
D7E117D8
18400001
D7E1F7F8
A84242C0
9FC00424
D7E14FFC
D7E177DC
D7E197E0
D7E1A7E4
D7E1B7E8
D7E1C7EC
D7E1D7F0
D7E1E7F4
84620000
A8BE0000
D7E10FD4
9C800000
9C21FFD4
07FFEE67
1B400001
84C20000
1B800001
9C860354
9C6603BC
9CA602EC
AB5A1D9C
9F00330E
9EC0ABCD
9E801234
9E40E66D
9DC0DEEC
AB9C4B80
D4062008
D406180C
9C80000B
9C600005
D4062804
D406D034
DC06C0AC
DC06B0AE
DC06A0B0
DC0690B2
DC0670B4
DC0618B6
DC0620B8
847C0000
A8BE0000
9CE00000
9D000001
D40638A4
D40640A8
07FFEE46
9C800000
847C0000
84420000
9C8303BC
9D000005
D403200C
9C80000B
DC0340B6
DC0320B8
18800001
9CC302EC
A8845130
9CA30354
D4041000
18800001
9CE00000
A884512C
9D000001
DC03C0AC
DC03B0AE
DC03A0B0
DC0390B2
DC0370B4
D40338A4
D40340A8
D403D034
D4041000
D4033004
D4032808
9C21002C
8521FFFC
8421FFD4
8441FFD8
85C1FFDC
8641FFE0
8681FFE4
86C1FFE8
8701FFEC
8741FFF0
8781FFF4
44004800
87C1FFF8
18600001
D7E10FFC
A863512C
9C21FFFC
85630000
9C210004
44004800
8421FFFC
D7E10FFC
9C21FFFC
9C210004
44004800
8421FFFC
D7E14FFC
D7E117F8
D7E10FF4
9C21FFF4
07FFFFF7
9C400000
18800000
18600001
A884FF30
A8635148
D4032018
18600001
A8635134
D4031000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E14FFC
D7E117F8
D7E10FF4
07FFFEFF
9C21FFF4
040000CB
A84B0000
9C21000C
E0421000
8521FFFC
8421FFF4
E1625804
44004800
8441FFF8
D7E14FFC
D7E117F8
D7E10FF4
A8430000
9C21FFF4
040000CB
A4630001
B8620041
07FFFEFA
A4630001
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
44004800
E1600004
44004800
E1600004
44004800
A9600001
44004800
85630000
44004800
D4032000
85630000
E40B2000
0C000003
15000000
D4032800
44004800
15000000
E0800004
03FFFFF8
9CA00001
9C63FFFE
D7E117FC
18400001
B8630002
A8425148
D7E10FF8
E0631000
9C21FFF8
D4032000
9C210008
8421FFF8
44004800
8441FFFC
18A00001
D7E10FF8
A8A55120
D7E117FC
84650000
9C21FFF8
9C630001
9C805000
D4051800
B4640000
18402FFF
A842FFFF
E0631003
18406000
E0631004
C0041800
9C210008
8421FFF8
44004800
8441FFFC
D7E197F8
D7E14FFC
D7E10FEC
D7E117F0
D7E177F4
9E400001
9C21FFEC
B4B20000
B8A5004A
E0A59003
BC050000
10000020
18400001
A8830000
A842070C
19C00001
84620000
07FFD19F
18400FFF
A842FFFF
A9CE5120
E16B1003
9C405000
D40E5804
C0025800
18800001
9C400000
9C600005
A88403A0
D40E1000
07FFFFC1
15000000
9C605001
D40E9008
C0031000
A9620000
9C210014
8521FFFC
8421FFEC
8441FFF0
85C1FFF4
44004800
8641FFF8
03FFFFF9
9D60FFFF
A8830000
18600001
D7E117F8
A863070C
18400FFF
D7E14FFC
D7E10FF4
84630000
9C21FFF4
07FFD17A
A842FFFF
9C805000
E16B1003
B4640000
1840F000
E0631003
E0635804
C0041800
18600001
A8635120
D4035804
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E14FFC
D7E10FF8
A8830000
9C21FFF8
07FFFF94
9C600005
9C210008
8521FFFC
44004800
8421FFF8
18800001
D7E10FF8
A8845120
D7E117FC
9CA05000
9C21FFF8
D4041808
B4850000
B8C4005E
BC060000
10000007
B863001E
18403FFF
A842FFFF
E0841003
E0641804
C0051800
9C210008
8421FFF8
44004800
8441FFFC
D7E10FF8
D7E117FC
9CA05000
9C21FFF8
B4650000
18403FFF
A842FFFF
E0831003
18600001
18402000
A8635120
84630008
B863001E
E0631004
E0632004
C0051800
9C800011
B4640000
A8630002
C0041800
9C210008
8421FFF8
44004800
8441FFFC
D7E10FF8
D7E117FC
9C600011
9C21FFF8
B5630000
9C40FFFD
E08B1003
C0032000
9C210008
B96B0041
8421FFF8
A56B0001
44004800
8441FFFC
D7E10FFC
9C800011
9C21FFFC
B4640000
A8630002
C0041800
9C210004
44004800
8421FFFC
D7E10FF8
D7E117FC
9C805000
9C21FFF8
B4640000
18403FFF
A842FFFF
E0631003
C0041800
9C210008
8421FFF8
44004800
8441FFFC
D7E10FF8
D7E117FC
9C805000
9C21FFF8
B4640000
1840EFFF
A842FFFF
E0631003
C0041800
9C800000
9C605001
C0032000
9C210008
8421FFF8
44004800
8441FFFC
18600001
D7E10FFC
A8635120
9C21FFFC
85630000
9C210004
44004800
8421FFFC
18600001
D7E117FC
A8635120
9C400000
D7E10FF8
9C21FFF8
D4031000
9C210008
8421FFF8
44004800
8441FFFC
04000000
02FAF080
90000000
0001C200
00000002
1500000C
15000000
44004800
15000000
44004800
15000000
D7E14FFC
D7E10FF8
07FFE882
9C21FFF8
9C210008
8521FFFC
44004800
8421FFF8
9C21FFF8
D4014800
D4017004
9CA30000
9DC00000
E5850000
0C000004
9C600000
9DC00001
E0A02802
E5840000
0C000004
15000000
9DCE0001
E0802002
07FFD0C7
9C650000
BC0E0001
0C000003
15000000
E1605802
85210000
85C10004
44004800
9C210008
9C21FFF8
D4014800
D4017004
9DC00000
E5830000
0C000004
15000000
9DC00001
E0601802
E5840000
0C000003
15000000
E0802002
07FFD0B0
15000000
BC0E0001
0C000003
9D670000
E1605802
85210000
85C10004
44004800
9C210008
D7E117EC
1840000F
D7E197F4
A842FFFF
BA43005F
E0E31003
E1651003
B9A5005F
B9870003
B9E6005D
B8630054
B8E4005D
B8A50054
B96B0003
D7E177F0
D7E14FFC
D7E10FE8
D7E1A7F8
E4326800
9C21FFE8
A44307FF
A9120000
E0EC3804
B9C40003
A4A507FF
E16B7804
0C000099
B8C60003
E0622802
BDA30000
100000F8
BC250000
1000003C
BC0207FF
E08B3004
BC040000
0C0000C6
9C63FFFF
A46E0007
BC230000
0C000088
18800080
A46E000F
BC230004
0C0000E7
18A00080
9C8E0004
E4847000
0C0000B8
9C600001
E0E71800
18A00080
A9120000
E0672803
A9C40000
BC030000
1000006E
B887001D
9C420001
BC0207FF
100000F3
1860FF7F
B9CE0043
A863FFFF
A44207FF
E0E71803
B887001D
B8E70043
E1C47004
1880000F
A884FFFF
E0E72003
A46207FF
1840000F
B8630014
A842FFFF
B908001F
E0E71003
9C210018
E0471804
A8AE0000
E0424004
8521FFFC
A8820000
8421FFE8
E1640004
E1850004
8441FFEC
85C1FFF0
8641FFF4
44004800
8681FFF8
13FFFFCA
BD430038
19000080
E16B4004
100000E3
BD43001F
1000010F
9C83FFE0
9D000020
E0861848
E1081802
E06B1848
E0A64008
E16B4008
E0C02802
E16B2004
E0A62804
B8A5005F
E08B2804
E08E2002
E0E71802
E4447000
10000003
9C600001
9C600000
E0E71802
A9C40000
18800080
E0672003
BC030000
10000091
A46E0007
18A0007F
A8A5FFFF
E2872803
BC140000
100000B2
15000000
07FFD063
A8740000
9C6BFFF8
BD43001F
100000B3
9C800028
E2941808
E1645802
E5421800
E16E5848
E1CE1808
100000B1
E16BA004
E0431002
9CE20001
BD47001F
100000D1
9C82FFE1
9C60001F
E0AE3848
E0431002
E0EB3848
E08E1008
E16B1008
9C400000
E1C02002
E1655804
E1CE2004
E1CE1848
03FFFF87
E1CB7004
18E0007F
9DC0FFF8
A8E7FFFF
9C4007FF
B887001D
B9CE0043
BC0207FF
B8E70043
10000036
E1C47004
1860000F
A44207FF
A863FFFF
03FFFF9A
E0E71803
A9120000
03FFFF86
E0672003
E0822802
BDA40000
10000094
BC250000
0C00003E
E06B3004
BC0207FF
13FFFF6C
18600080
E16B1804
BD440038
0C0000EA
BD44001F
E0CB3004
9C800000
E0603002
E0C33004
B866005F
E0637000
E0E43800
E4837000
10000003
9C800001
9C800000
E0E72000
A9C30000
18800080
E0672003
BC030000
1000003B
A46E0007
9C420001
BC0207FF
10000157
18A0FF7F
A46E0001
A8A5FFFF
E0E72803
B8AE0041
B887001F
B8E70041
E1C51804
03FFFF49
E1CE2004
E06E3804
BC030000
100001AD
18800008
18A0000F
E0E72004
A8A5FFFF
03FFFF62
E0E72803
03FFFF4A
9C600000
BC230000
10000074
BC0207FF
E0CE3002
E0E75802
E4467000
0C0000C6
9CA00001
E0E72802
03FFFF84
A9C60000
BC030000
13FFFF30
9C84FFFF
BC240000
100000D1
BC0207FF
E0C67000
E0EB3800
E4867000
10000003
9CA00001
A8A40000
E0E72800
03FFFFCB
A9C60000
E0E32004
BC070000
100001D4
15000000
A8E30000
A9C40000
A46E0007
BC230000
0FFFFF99
A9120000
A46E000F
BC230004
13FFFF1F
9C8E0004
18A00080
A9120000
03FFFF23
E0672803
BC030000
0C000067
9C820001
A48407FF
BD440001
0C0000D2
E08E3002
E2875802
E4447000
10000003
9CA00001
A8A30000
E2942802
19000080
E0744003
BC030000
1000007A
E16B3802
E1C67002
E44E3000
0C00009E
9C800001
E28B2002
03FFFF52
AA4D0000
9CE00000
03FFFF18
A9C70000
07FFCFB3
A86E0000
9D6B0020
9C6BFFF8
BD43001F
0FFFFF51
9C800028
9D6BFFD8
E5421800
E16E5808
0FFFFF53
9DC00000
1900FF7F
E0421802
A908FFFF
03FFFEE5
E0EB4003
E0CB3004
9C600000
E0803002
E0C43004
03FFFF28
B886005F
BC040000
0C0000C3
BC220000
9CA20001
A46507FF
BD430001
0C000083
BC0507FF
100000E3
E0C67000
E0EB3800
E4867000
10000003
9C400001
A8440000
E0E71000
B8C60041
B9C7001F
A8450000
B8E70041
03FFFEC9
E1CE3004
0FFFFF01
BD430038
03FFFEC6
A46E0007
BC070020
1000006A
E08B2048
9C60003F
E0431002
E16B1008
E1CB7004
9CE00000
E0607002
A8470000
E1C37004
B9CE005F
03FFFF9B
E1CE2004
BC030020
1000005E
E0AB2048
9C800040
E0641802
E16B1808
E0CB3004
9C600000
E0803002
E0C43004
B886005F
03FFFEF3
E0842804
BC220000
0C000039
E0477004
BC0507FF
10000086
E0601802
18400080
E0E71004
BD430038
100000A7
BD43001F
10000124
9C43FFE0
9C800020
E10E1848
E0841802
E0671848
E04E2008
E0872008
E0E01002
E0844004
E0471004
B842005F
E1C41004
E1C67002
E06B1802
E44E3000
10000003
9CE00001
9CE00000
E0E33802
A8450000
03FFFED9
AA4D0000
E0F42004
BC070000
0FFFFEDD
A9C40000
A9070000
A9C70000
03FFFEFF
A8470000
10000051
BC040020
9CA00020
E0662048
E0A52002
E08B2048
E0C62808
E16B2808
E0A03002
E06B1804
E0C53004
B8C6005F
03FFFF11
E0633004
03FFFF3C
A8A30000
BC020000
1000004F
AC63FFFF
BC230000
1000004A
BC0507FF
E1C67002
E0EB3802
E44E3000
10000003
9C400001
A8430000
E0E71002
AA4D0000
03FFFEB1
A8450000
03FFFF64
9C800000
0FFFFEF4
BD440038
03FFFE5B
A46E0007
03FFFF9B
9D600000
03FFFFA7
9D600000
BC220000
100000BE
E0677004
BC030000
100000EE
E06B3004
BC030000
13FFFE4E
A46E0007
E0A67000
E0EB3800
E4857000
10000003
9C800001
A8820000
E0E72000
18800080
E0672003
BC030000
100000F8
15000000
1900FF7F
A9C50000
A908FFFF
9C400001
03FFFE3B
E0E74003
BC220000
10000031
E0677004
BC230000
10000064
E06B3004
BC030000
100000C6
AA4D0000
A8EB0000
03FFFE2F
A9C60000
9C64FFE0
100000B1
E0AB1848
9C600040
E0832002
E16B2008
E0CB3004
9C800000
E0603002
E0C33004
B866005F
03FFFEC1
E0632804
0FFFFF81
BD430038
A8EB0000
A9C60000
A8450000
03FFFE1B
AA4D0000
1000002B
BC0507FF
E0477004
BC020000
10000079
AC84FFFF
BC240000
10000074
BC0507FF
E1CE3000
E0EB3800
E48E3000
10000003
9C400001
A8440000
E0E71000
03FFFEB0
A8450000
E0477004
BC220000
1000004B
E06B3004
E10B3004
BC080000
13FFFE7C
A8EB0000
A9C60000
AA4D0000
03FFFDFD
9C4007FF
9CE00000
03FFFE79
A9C70000
E0E77004
9C600000
E1C03802
E1CE3804
03FFFF64
B9CE005F
A8E40000
A8450000
03FFFE6F
A9C40000
10000052
E0802002
18400080
E0E71004
BD440038
10000081
BD44001F
1000008C
9C44FFE0
9C600020
E18E2048
E0632002
E0872048
E04E1808
E0671808
E0E01002
E0636004
E0471004
B842005F
E1C31004
E1CE3000
E1645800
E48E3000
10000003
9CE00001
9CE00000
E0EB3800
03FFFE7A
A8450000
BC030000
13FFFDD1
A46E0007
E08E3002
E0675802
E4447000
10000003
9CA00001
A8A20000
E0632802
19000080
E0A34003
BC050000
13FFFEA2
E1C67002
E0EB3802
E44E3000
10000003
9C800001
9C800000
E0E72002
03FFFDBC
AA4D0000
BC030000
13FFFDB9
9C4007FF
B8470043
18800008
B9CE0043
E0622003
B8E7001D
BC030000
1000000D
E1C77004
B88B0043
18A00008
E0642803
BC230000
10000008
B8620003
B8C60043
B96B001D
A8440000
AA4D0000
E1CB3004
B8620003
B8EE005D
9C4007FF
B9CE0003
03FFFDA0
E0E71804
0FFFFFB5
BD440038
A8EB0000
A9C60000
03FFFD9A
A8450000
A8E30000
03FFFDB9
A9C30000
E0477004
BC020000
10000034
E06B3004
BC030000
13FFFD90
9C4007FF
B8470043
18800008
B9CE0043
E0622003
B8E7001D
BC030000
13FFFFE4
E1C77004
B88B0043
18A00008
E0642803
BC230000
13FFFFDF
B8620003
B8C60043
B96B001D
A8440000
03FFFFD9
E1CB3004
03FFFF54
9D600000
BC030020
1000002A
E0471048
9C800040
E0641802
E0E71808
E1C77004
9C600000
E0807002
E1C47004
B9CE005F
03FFFEDE
E1CE1004
A9020000
A8E20000
03FFFDE9
A9C20000
E0E77004
9C800000
E1C03802
E1CE3804
03FFFF8A
B9CE005F
A8EB0000
03FFFD61
A9C60000
A8EB0000
A9C60000
03FFFD5D
9C4007FF
BC040020
10000013
E0471048
9C600040
E0832002
E0E72008
E1C77004
9C800000
E0607002
E1C37004
B9CE005F
03FFFF76
E1CE1004
03FFFFDB
9CE00000
A9070000
03FFFDCA
A9C70000
03FFFE2D
A9C50000
03FFFFF2
9CE00000
D7E117FC
1840000F
B8E30054
A842FFFF
B9050054
E1831003
A4E707FF
1840000F
D7E10FF8
A842FFFF
BC2707FF
E1A51003
9C21FFF8
B863005F
A50807FF
0C00000C
B8A5005F
BC2807FF
0C000011
E1ED3004
E4274000
0C000014
9D600001
9C210008
8421FFF8
44004800
8441FFFC
E1EC2004
BC2F0000
13FFFFFA
9D600001
BC2807FF
13FFFFF5
E4274000
E1ED3004
BC2F0000
13FFFFF3
9D600001
E4274000
13FFFFF0
15000000
E42C6800
10000011
E0C62005
E1003002
E0C83004
B8C6005F
BC260000
1000000B
E4032800
1000000E
BC270000
13FFFFE3
15000000
E08C2004
E1602002
E08B2004
03FFFFDE
B964005F
9C210008
9D600001
8421FFF8
44004800
8441FFFC
03FFFFD7
A9660000
D7E117FC
1840000F
B9030054
A842FFFF
B9650054
E1A31003
A50807FF
1840000F
D7E10FF8
A842FFFF
BC2807FF
E1851003
9C21FFF8
B863005F
A56B07FF
0C000018
B8A5005F
BC2B07FF
0C000033
BC280000
10000019
BC2B0000
E0ED2004
BC2B0000
E1E03802
E0EF3804
ACE7FFFF
10000020
B8E7005F
E1EC3004
BC2F0000
1000001D
BC270000
0C000013
BC030000
9C210008
8421FFF8
44004800
8441FFFC
E0ED2004
BC270000
1000004E
BC0B07FF
1000001A
BC2B0000
1000001F
E4032800
E0EC3004
BC070000
0C00001B
E4032800
BC030000
13FFFFEF
9D600001
9C210008
9D60FFFF
8421FFF8
44004800
8441FFFC
BC270000
0C00000F
BC050000
13FFFFE5
9D60FFFF
9C210008
9D600001
8421FFF8
44004800
8441FFFC
E0EC3004
BC270000
10000030
BC080000
13FFFFCE
E0ED2004
E4032800
0FFFFFE8
BC030000
E5A85800
0FFFFFE5
BC030000
E5685800
0C000021
BC030000
E44D6000
13FFFFDF
BC030000
E0AD6005
E0E02802
E0A72804
ACA5FFFF
B8A5005F
BC050000
10000009
E4443000
10000003
9CE00001
9CE00000
A4E700FF
BC070000
0FFFFFD0
BC030000
E48D6000
1000000C
BC030000
BC050000
1000000F
E4462000
10000003
9C800001
9C800000
A48400FF
BC040000
10000008
BC030000
13FFFFB0
9D60FFFF
03FFFFCC
9C210008
03FFFFAC
9D60FFFE
03FFFFAA
9D600000
D7E117FC
1840000F
B9030054
A842FFFF
B8E50054
E1A31003
A50807FF
1840000F
D7E10FF8
A842FFFF
BC2807FF
E1851003
9C21FFF8
B863005F
A4E707FF
0C000017
B8A5005F
BC2707FF
0C000033
BC280000
10000019
BC270000
E16D2004
BC270000
E1E05802
E16F5804
AD6BFFFF
0C000020
B96B005F
BC2B0000
0C000015
BC050000
0C000054
9D60FFFF
9C210008
8421FFF8
44004800
8441FFFC
E1ED2004
BC2F0000
13FFFFFA
9D600002
BC0707FF
1000001A
BC270000
10000007
E4032800
E16C3004
BC0B0000
10000006
BC030000
E4032800
1000001A
E5A83800
BC030000
13FFFFEB
9D600001
03FFFFE9
9D60FFFF
E1EC3004
BC2F0000
13FFFFE1
BC2B0000
0FFFFFF7
A9670000
9C210008
8421FFF8
44004800
8441FFFC
E1EC3004
BC2F0000
13FFFFDB
9D600002
BC080000
13FFFFCC
E4032800
03FFFFE8
15000000
0FFFFFE9
BC030000
E5683800
0C000021
BC030000
E44D6000
13FFFFE3
BC030000
E0AD6005
E0E02802
E0A72804
ACA5FFFF
B8A5005F
BC050000
10000009
E4443000
10000003
9CE00001
9CE00000
A4E700FF
BC070000
0FFFFFD4
BC030000
E48D6000
1000000C
BC030000
BC050000
1000000D
E4462000
10000003
9C800001
9C800000
A48400FF
BC040000
10000006
BC030000
13FFFFB0
9D60FFFF
03FFFFAE
9D600001
03FFFFAC
9D600000
B8A30054
D7E117FC
1840000F
A4A507FF
D7E10FF8
A842FFFF
BDA503FE
E0C31003
9C21FFF8
B863005F
10000010
9D600000
BDA5041D
0C000011
9CE00433
18400010
E0E72802
BD47001F
0C000013
E0C61004
9D600413
E16B2802
E1665848
E0C01802
E16B3005
E16B1800
9C210008
8421FFF8
44004800
8441FFFC
9C210008
18407FFF
8421FFF8
A842FFFF
E1631000
44004800
8441FFFC
9CA5FBED
E1643848
E0A62808
03FFFFEF
E16B2804
D7E117F4
D7E14FFC
D7E10FF0
D7E177F8
BC030000
9C21FFF0
10000018
A8430000
B9C3005F
BC0E0000
10000003
15000000
E0401802
07FFCC98
A8620000
9C60041E
BD4B000A
10000021
E0635802
9CA0000B
9C8B0015
E1655802
18A0000F
E1625848
A8A5FFFF
E0822008
A46307FF
A84E0000
00000004
E16B2803
A9620000
A8820000
18A0000F
A46307FF
A8A5FFFF
B8630014
E16B2803
B842001F
E06B1804
9C210010
E0431004
A8E40000
A8C20000
8521FFFC
8421FFF0
E1660004
E1870004
8441FFF4
44004800
85C1FFF8
9D6BFFF5
18A0000F
E1625808
A8A5FFFF
A46307FF
A84E0000
9C800000
03FFFFE7
E16B2803
D7E117F8
18400001
D7E14FFC
A8424294
D7E10FF4
8462FFFC
9C21FFF4
BC23FFFF
0C000008
9C42FFFC
48001800
9C42FFFC
84620000
BC23FFFF
13FFFFFC
15000000
9C21000C
8521FFFC
8421FFF4
44004800
8441FFF8
D7E14FFC
D7E10FF8
9C21FFF8
9C210008
8521FFFC
44004800
8421FFF8
9C21FFFC
D4014800
07FFC1E3
15000000
85210000
44004800
9C210004
57726974
65333220
61646472
6573733A
20253038
780A0052
65616433
32206164
64726573
733A2025
3038780A
00496E63
6F727265
63742076
616C7565
20253038
78206174
20616464
72657373
20253038
782C2065
78706563
74656420
25303878
0A005772
69746531
36206164
64726573
733A2025
3038780A
00526561
64313620
61646472
6573733A
20253038
780A0049
6E636F72
72656374
2076616C
75652025
30347820
61742061
64647265
73732025
3038782C
20657870
65637465
64202530
34780A00
57726974
65382061
64647265
73733A20
25303878
0A005265
61643820
61646472
6573733A
20253038
780A0049
6E636F72
72656374
2076616C
75652025
30327820
61742061
64647265
73732025
3038782C
20657870
65637465
64202530
32780A00
41646472
6573733A
20253038
780A0044
69652074
656D7065
72617475
72653A20
25662043
64656720
28726177
2076616C
75653A20
25303878
290A0000
407F7F99
9999999A
40F00000
40711266
66666666
48656C6C
6F20576F
726C6421
00002DD8
00002D10
00002D98
00002BD4
00002D98
00002D80
00002D98
00002BD4
00002D10
00002D10
00002D80
00002BD4
00002BE4
00002BE4
00002BE4
00002DA8
0000397C
00003968
00003968
00003954
00003798
00003798
0000393C
00003954
00003798
0000393C
00003798
00003954
0000379C
0000379C
0000379C
00003C10
00010202
03030303
04040404
04040404
05050505
05050505
05050505
05050505
06060606
06060606
06060606
06060606
06060606
06060606
06060606
06060606
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
000142C4
43000A00
494E4600
696E6600
4E414E00
6E616E00
30313233
34353637
38394142
43444546
00303132
33343536
37383961
62636465
6600286E
756C6C29
00300000
00005504
00005980
00005980
00005518
00005980
00005980
00005980
00005980
00005980
00005980
00005160
000052A0
00005980
00005190
00005524
00005980
00005580
00005600
00005600
00005600
00005600
00005600
00005600
00005600
00005600
00005600
00005980
00005980
00005980
00005980
00005980
00005980
00005980
00005980
00005980
00005980
00005640
00005688
00005980
00005688
00005980
00005980
00005980
00005980
00005764
00005980
00005980
00005770
00005980
00005980
00005980
00005980
00005980
000057B0
00005980
00005980
000057F4
00005980
00005980
00005980
00005980
00005980
00005980
00005980
00005980
00005980
00005980
00005860
000058A8
00005688
00005688
00005688
000058E8
000058A8
00005980
00005980
00005154
00005980
00005940
0000558C
000055BC
00005154
00005980
000052AC
00005980
0000543C
00005980
00005980
000058F4
30303030
30303030
30303030
30303030
20202020
20202020
20202020
20202020
496E6669
6E697479
004E614E
3FF80000
3FD287A7
636F4361
3FC68A28
8B60C8B3
3FD34413
509F79FB
3FF00000
40240000
401C0000
40140000
3FE00000
7FFFFFFF
504F5349
58002E00
3FF00000
40240000
00000005
00000019
0000007D
3C9CD2B2
97D889BC
3949F623
D5A8A733
32A50FFD
44F4A73D
255BBA08
CF8C979D
0AC80628
64AC6F43
4341C379
37E08000
4693B8B5
B5056E17
4D384F03
E93FF9F5
5A827748
F9301D32
75154FDD
7F73BF3C
3FF00000
40240000
40590000
408F4000
40C38800
40F86A00
412E8480
416312D0
4197D784
41CDCD65
4202A05F
20000000
42374876
E8000000
426D1A94
A2000000
42A2309C
E5400000
42D6BCC4
1E900000
430C6BF5
26340000
4341C379
37E08000
43763457
85D8A000
43ABC16D
674EC800
43E158E4
60913D00
4415AF1D
78B58C40
444B1AE4
D6E2EF50
4480F0CF
064DD592
44B52D02
C7E14AF6
44EA7843
79D99DB4
0000E71C
0000E938
0000E938
0000E778
0000E938
0000E938
0000E938
0000E938
0000E938
0000E938
0000E580
0000E5B8
0000E938
0000E5AC
0000E784
0000E938
0000E730
0000E5C4
0000E5C4
0000E5C4
0000E5C4
0000E5C4
0000E5C4
0000E5C4
0000E5C4
0000E5C4
0000E938
0000E938
0000E938
0000E938
0000E938
0000E938
0000E938
0000E938
0000E938
0000E938
0000E60C
0000E938
0000E938
0000E938
0000E938
0000E938
0000E938
0000E938
0000E938
0000E938
0000E938
0000DD4C
0000E938
0000E938
0000E938
0000E938
0000E938
0000DD10
0000E938
0000E938
0000E650
0000E938
0000E938
0000E938
0000E938
0000E938
0000E938
0000E938
0000E938
0000E938
0000E938
0000E6AC
0000E6E4
0000E938
0000E938
0000E938
0000E818
0000E6E4
0000E938
0000E938
0000DD04
0000E938
0000E86C
0000DD50
0000E7E0
0000DD04
0000E938
0000E898
0000E938
0000DD14
0000E938
0000E938
0000E824
30303030
30303030
30303030
30303030
20202020
20202020
20202020
20202020
FFFFFFFF
FFFFFFFF
00002000
00002000
3F065B4F
666D7D07
7F6F777C
395E7971
000142C4
000145B0
00014618
00014680
00011D9C
00000001
330EABCD
1234E66D
DEEC0005
000B0000
41534349
49000000
41534349
49000000
00011FD2
00011D9F
00011D9F
00011D9F
00011D9F
00011D9F
00011D9F
00011D9F
00011D9F
00011D9F
7F7F7F7F
7F7F7F7F
7F7F7F7F
7F7F0000
00000001
FFFFFFFF
00020000
0001476C
0001476C
00014774
00014774
0001477C
0001477C
00014784
00014784
0001478C
0001478C
00014794
00014794
0001479C
0001479C
000147A4
000147A4
000147AC
000147AC
000147B4
000147B4
000147BC
000147BC
000147C4
000147C4
000147CC
000147CC
000147D4
000147D4
000147DC
000147DC
000147E4
000147E4
000147EC
000147EC
000147F4
000147F4
000147FC
000147FC
00014804
00014804
0001480C
0001480C
00014814
00014814
0001481C
0001481C
00014824
00014824
0001482C
0001482C
00014834
00014834
0001483C
0001483C
00014844
00014844
0001484C
0001484C
00014854
00014854
0001485C
0001485C
00014864
00014864
0001486C
0001486C
00014874
00014874
0001487C
0001487C
00014884
00014884
0001488C
0001488C
00014894
00014894
0001489C
0001489C
000148A4
000148A4
000148AC
000148AC
000148B4
000148B4
000148BC
000148BC
000148C4
000148C4
000148CC
000148CC
000148D4
000148D4
000148DC
000148DC
000148E4
000148E4
000148EC
000148EC
000148F4
000148F4
000148FC
000148FC
00014904
00014904
0001490C
0001490C
00014914
00014914
0001491C
0001491C
00014924
00014924
0001492C
0001492C
00014934
00014934
0001493C
0001493C
00014944
00014944
0001494C
0001494C
00014954
00014954
0001495C
0001495C
00014964
00014964
0001496C
0001496C
00014974
00014974
0001497C
0001497C
00014984
00014984
0001498C
0001498C
00014994
00014994
0001499C
0001499C
000149A4
000149A4
000149AC
000149AC
000149B4
000149B4
000149BC
000149BC
000149C4
000149C4
000149CC
000149CC
000149D4
000149D4
000149DC
000149DC
000149E4
000149E4
000149EC
000149EC
000149F4
000149F4
000149FC
000149FC
00014A04
00014A04
00014A0C
00014A0C
00014A14
00014A14
00014A1C
00014A1C
00014A24
00014A24
00014A2C
00014A2C
00014A34
00014A34
00014A3C
00014A3C
00014A44
00014A44
00014A4C
00014A4C
00014A54
00014A54
00014A5C
00014A5C
00014A64
00014A64
00014A6C
00014A6C
00014A74
00014A74
00014A7C
00014A7C
00014A84
00014A84
00014A8C
00014A8C
00014A94
00014A94
00014A9C
00014A9C
00014AA4
00014AA4
00014AAC
00014AAC
00014AB4
00014AB4
00014ABC
00014ABC
00014AC4
00014AC4
00014ACC
00014ACC
00014AD4
00014AD4
00014ADC
00014ADC
00014AE4
00014AE4
00014AEC
00014AEC
00014AF4
00014AF4
00014AFC
00014AFC
00014B04
00014B04
00014B0C
00014B0C
00014B14
00014B14
00014B1C
00014B1C
00014B24
00014B24
00014B2C
00014B2C
00014B34
00014B34
00014B3C
00014B3C
00014B44
00014B44
00014B4C
00014B4C
00014B54
00014B54
00014B5C
00014B5C
00014B64
00014B64
0000F5D0
00015008
000151C0
00014B84
00014E70
00014ED8
00014F40
00011D9C
00000001
330EABCD
1234E66D
DEEC0005
000B0000
	 
