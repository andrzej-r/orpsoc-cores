@00000000
18000000
18200000
18400000
18600000
18800000
18A00000
18C00000
A8C60100
44003000
15000000
	 
