@00000000
18000000
18A00000
A8A50800
18800000
C0802002
9C840010
E4842800
13FFFFFD
15000000
B4800011
A8840010
C0002011
B4800011
A8840008
C0002011
18A00000
A8A50800
18800000
C0602003
9C840010
E4842800
13FFFFFD
15000000
18200000
A821025C
18400000
A8420300
18600800
A8630000
18A0FFFF
A8A5FFFF
18C09100
A8C62000
D4062804
18E09200
A8E70000
18A00000
A8A50001
D4072800
D4021000
A4A2FFFF
E4050000
0C000004
15000000
0400000A
15000000
9C420004
E4021800
0FFFFFF7
15000000
04000004
15000000
04000000
15000000
E1890004
B8820040
04000019
9CA7003C
B8820044
04000016
9CA70038
B8820048
04000013
9CA70034
B882004C
04000010
9CA70030
B8820050
0400000D
9CA7002C
B8820054
0400000A
9CA70028
B8820058
04000007
9CA70024
B882005C
04000004
9CA70020
44006000
15000000
A484000F
E0840800
8C840000
D4052000
44004800
15000000
3F065B4F
666D7D07
7F6F777C
395E7971
	 
