@00000000
18000000
1880DEAD
A884BEEF
15000000
D4002000
D4002004
D4002008
D400200C
D4002010
D4002014
D4002018
D400201C
D4002020
D4002024
D4002028
D400202C
84600000
84600004
84600008
8460000C
84600040
84600044
84600048
8460004C
84600040
84600044
84600048
8460004C
84600000
84600004
84600008
8460000C
18A0F000
A8A50400
1880F000
C0802002
9C840010
E4842800
13FFFFFD
15000000
B4800011
A8840010
C0002011
B4800011
A8840008
C0002011
18A00000
A8A50200
18800000
C0602003
9C840010
E4842800
13FFFFFD
15000000
1880DEAD
A884BEEF
1880DEAD
A884BEEF
D4002000
D4002004
D4002008
D400200C
D4002010
D4002014
D4002018
D400201C
D4002020
D4002024
D4002028
D400202C
84600000
84600004
84600008
8460000C
84600040
84600044
84600048
8460004C
84600040
84600044
84600048
8460004C
84600000
84600004
84600008
8460000C
1880BEEF
A884DEAD
03FFFFE0
15000000
	 
